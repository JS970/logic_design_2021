// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Thu Nov 25 22:01:41 2021"

module six_bit_decoder(
	Din,
	D1,
	D16,
	D15,
	D14,
	D13,
	D12,
	D11,
	D10,
	D9,
	D8,
	D7,
	D6,
	D5,
	D4,
	D3,
	D2,
	D25,
	D33,
	D41,
	D49,
	D57,
	D17,
	D18,
	D19,
	D20,
	D21,
	D22,
	D23,
	D24,
	D26,
	D27,
	D28,
	D29,
	D30,
	D31,
	D32,
	D34,
	D35,
	D36,
	D37,
	D38,
	D39,
	D40,
	D42,
	D43,
	D44,
	D45,
	D46,
	D47,
	D48,
	D50,
	D51,
	D52,
	D53,
	D54,
	D55,
	D56,
	D58,
	D59,
	D60,
	D61,
	D62,
	D63,
	D64
);


input wire	[5:0] Din;
output wire	D1;
output wire	D16;
output wire	D15;
output wire	D14;
output wire	D13;
output wire	D12;
output wire	D11;
output wire	D10;
output wire	D9;
output wire	D8;
output wire	D7;
output wire	D6;
output wire	D5;
output wire	D4;
output wire	D3;
output wire	D2;
output wire	D25;
output wire	D33;
output wire	D41;
output wire	D49;
output wire	D57;
output wire	D17;
output wire	D18;
output wire	D19;
output wire	D20;
output wire	D21;
output wire	D22;
output wire	D23;
output wire	D24;
output wire	D26;
output wire	D27;
output wire	D28;
output wire	D29;
output wire	D30;
output wire	D31;
output wire	D32;
output wire	D34;
output wire	D35;
output wire	D36;
output wire	D37;
output wire	D38;
output wire	D39;
output wire	D40;
output wire	D42;
output wire	D43;
output wire	D44;
output wire	D45;
output wire	D46;
output wire	D47;
output wire	D48;
output wire	D50;
output wire	D51;
output wire	D52;
output wire	D53;
output wire	D54;
output wire	D55;
output wire	D56;
output wire	D58;
output wire	D59;
output wire	D60;
output wire	D61;
output wire	D62;
output wire	D63;
output wire	D64;

wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_131;





mux16bit	b2v_inst(
	.A(Din[0]),
	.B(Din[1]),
	.C(Din[2]),
	.D(Din[3]),
	.Q15(SYNTHESIZED_WIRE_21),
	.Q14(SYNTHESIZED_WIRE_23),
	.Q13(SYNTHESIZED_WIRE_5),
	.Q12(SYNTHESIZED_WIRE_7),
	.Q11(SYNTHESIZED_WIRE_9),
	.Q10(SYNTHESIZED_WIRE_11),
	.Q9(SYNTHESIZED_WIRE_13),
	.Q8(SYNTHESIZED_WIRE_15),
	.Q7(SYNTHESIZED_WIRE_17),
	.Q6(SYNTHESIZED_WIRE_19),
	.Q5(SYNTHESIZED_WIRE_99),
	.Q4(SYNTHESIZED_WIRE_117),
	.Q3(SYNTHESIZED_WIRE_127),
	.Q2(SYNTHESIZED_WIRE_129),
	.Q1(SYNTHESIZED_WIRE_1),
	.Q0(SYNTHESIZED_WIRE_3));

assign	D2 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_1;

assign	D1 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_3;

assign	D14 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_5;

assign	D13 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_7;

assign	D12 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_9;

assign	D11 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_11;

assign	D10 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_13;

assign	D9 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_15;

assign	D8 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_17;

assign	D7 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_19;

assign	D16 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_21;

assign	D15 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_23;

assign	SYNTHESIZED_WIRE_133 =  ~Din[4];

assign	SYNTHESIZED_WIRE_134 =  ~Din[5];

assign	SYNTHESIZED_WIRE_132 = SYNTHESIZED_WIRE_133 & SYNTHESIZED_WIRE_134;

assign	SYNTHESIZED_WIRE_137 = Din[4] & SYNTHESIZED_WIRE_134;

assign	SYNTHESIZED_WIRE_135 = SYNTHESIZED_WIRE_133 & Din[5];

assign	SYNTHESIZED_WIRE_136 = Din[4] & Din[5];

assign	D34 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_29;

assign	D33 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_31;

assign	D46 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_33;

assign	D45 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_35;

assign	D44 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_37;

assign	D43 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_39;

assign	D42 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_41;

assign	D41 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_43;

assign	D40 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_45;

assign	D39 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_47;

assign	D48 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_49;

assign	D47 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_51;

assign	D54 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_53;

assign	D53 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_55;

assign	D52 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_57;

assign	D51 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_59;

assign	D50 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_61;

assign	D49 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_63;

assign	D62 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_65;

assign	D61 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_67;

assign	D60 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_69;

assign	D59 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_71;


mux16bit	b2v_inst5(
	.A(Din[0]),
	.B(Din[1]),
	.C(Din[2]),
	.D(Din[3]),
	.Q15(SYNTHESIZED_WIRE_81),
	.Q14(SYNTHESIZED_WIRE_83),
	.Q13(SYNTHESIZED_WIRE_65),
	.Q12(SYNTHESIZED_WIRE_67),
	.Q11(SYNTHESIZED_WIRE_69),
	.Q10(SYNTHESIZED_WIRE_71),
	.Q9(SYNTHESIZED_WIRE_73),
	.Q8(SYNTHESIZED_WIRE_75),
	.Q7(SYNTHESIZED_WIRE_77),
	.Q6(SYNTHESIZED_WIRE_79),
	.Q5(SYNTHESIZED_WIRE_53),
	.Q4(SYNTHESIZED_WIRE_55),
	.Q3(SYNTHESIZED_WIRE_57),
	.Q2(SYNTHESIZED_WIRE_59),
	.Q1(SYNTHESIZED_WIRE_61),
	.Q0(SYNTHESIZED_WIRE_63));

assign	D58 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_73;

assign	D57 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_75;

assign	D56 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_77;

assign	D55 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_79;

assign	D64 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_81;

assign	D63 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_83;

assign	D22 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_85;

assign	D21 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_87;

assign	D20 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_89;

assign	D19 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_91;

assign	D38 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_93;

assign	D18 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_95;

assign	D17 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_97;

assign	D6 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_99;

assign	D30 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_101;

assign	D29 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_103;

assign	D28 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_105;

assign	D27 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_107;

assign	D26 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_109;

assign	D25 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_111;

assign	D24 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_113;

assign	D23 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_115;

assign	D5 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_117;

assign	D32 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_119;

assign	D31 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_121;


mux16bit	b2v_inst72(
	.A(Din[0]),
	.B(Din[1]),
	.C(Din[2]),
	.D(Din[3]),
	.Q15(SYNTHESIZED_WIRE_49),
	.Q14(SYNTHESIZED_WIRE_51),
	.Q13(SYNTHESIZED_WIRE_33),
	.Q12(SYNTHESIZED_WIRE_35),
	.Q11(SYNTHESIZED_WIRE_37),
	.Q10(SYNTHESIZED_WIRE_39),
	.Q9(SYNTHESIZED_WIRE_41),
	.Q8(SYNTHESIZED_WIRE_43),
	.Q7(SYNTHESIZED_WIRE_45),
	.Q6(SYNTHESIZED_WIRE_47),
	.Q5(SYNTHESIZED_WIRE_93),
	.Q4(SYNTHESIZED_WIRE_123),
	.Q3(SYNTHESIZED_WIRE_125),
	.Q2(SYNTHESIZED_WIRE_131),
	.Q1(SYNTHESIZED_WIRE_29),
	.Q0(SYNTHESIZED_WIRE_31));

assign	D37 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_123;


mux16bit	b2v_inst73(
	.A(Din[0]),
	.B(Din[1]),
	.C(Din[2]),
	.D(Din[3]),
	.Q15(SYNTHESIZED_WIRE_119),
	.Q14(SYNTHESIZED_WIRE_121),
	.Q13(SYNTHESIZED_WIRE_101),
	.Q12(SYNTHESIZED_WIRE_103),
	.Q11(SYNTHESIZED_WIRE_105),
	.Q10(SYNTHESIZED_WIRE_107),
	.Q9(SYNTHESIZED_WIRE_109),
	.Q8(SYNTHESIZED_WIRE_111),
	.Q7(SYNTHESIZED_WIRE_113),
	.Q6(SYNTHESIZED_WIRE_115),
	.Q5(SYNTHESIZED_WIRE_85),
	.Q4(SYNTHESIZED_WIRE_87),
	.Q3(SYNTHESIZED_WIRE_89),
	.Q2(SYNTHESIZED_WIRE_91),
	.Q1(SYNTHESIZED_WIRE_95),
	.Q0(SYNTHESIZED_WIRE_97));

assign	D36 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_125;

assign	D4 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_127;

assign	D3 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_129;

assign	D35 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_131;


endmodule
