// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Nov 24 20:57:16 2021"

module P(
	pin1,
	pin2,
	pin3,
	pin4,
	pin5,
	pin6,
	pin7,
	pin8,
	pin9,
	pin10,
	pin11,
	pin12,
	pin13,
	pin14,
	pin15,
	pin16,
	pin17,
	pin18,
	pin19,
	pin20,
	pin21,
	pin22,
	pin23,
	pin24,
	pin25,
	pin26,
	pin27,
	pin28,
	pin29,
	pin30,
	pin31,
	pin32,
	pout1,
	pout2,
	pout3,
	pout4,
	pout5,
	pout6,
	pout7,
	pout8,
	pout9,
	pout10,
	pout11,
	pout12,
	pout13,
	pout14,
	pout15,
	pout16,
	pout17,
	pout18,
	pout19,
	pout20,
	pout21,
	pout22,
	pout23,
	pout24,
	pout25,
	pout26,
	pout27,
	pout28,
	pout29,
	pout30,
	pout31,
	pout32
);


input wire	pin1;
input wire	pin2;
input wire	pin3;
input wire	pin4;
input wire	pin5;
input wire	pin6;
input wire	pin7;
input wire	pin8;
input wire	pin9;
input wire	pin10;
input wire	pin11;
input wire	pin12;
input wire	pin13;
input wire	pin14;
input wire	pin15;
input wire	pin16;
input wire	pin17;
input wire	pin18;
input wire	pin19;
input wire	pin20;
input wire	pin21;
input wire	pin22;
input wire	pin23;
input wire	pin24;
input wire	pin25;
input wire	pin26;
input wire	pin27;
input wire	pin28;
input wire	pin29;
input wire	pin30;
input wire	pin31;
input wire	pin32;
output wire	pout1;
output wire	pout2;
output wire	pout3;
output wire	pout4;
output wire	pout5;
output wire	pout6;
output wire	pout7;
output wire	pout8;
output wire	pout9;
output wire	pout10;
output wire	pout11;
output wire	pout12;
output wire	pout13;
output wire	pout14;
output wire	pout15;
output wire	pout16;
output wire	pout17;
output wire	pout18;
output wire	pout19;
output wire	pout20;
output wire	pout21;
output wire	pout22;
output wire	pout23;
output wire	pout24;
output wire	pout25;
output wire	pout26;
output wire	pout27;
output wire	pout28;
output wire	pout29;
output wire	pout30;
output wire	pout31;
output wire	pout32;


assign	pout1 = pin16;
assign	pout2 = pin7;
assign	pout3 = pin20;
assign	pout4 = pin21;
assign	pout5 = pin29;
assign	pout6 = pin12;
assign	pout7 = pin28;
assign	pout8 = pin17;
assign	pout9 = pin1;
assign	pout10 = pin15;
assign	pout11 = pin23;
assign	pout12 = pin26;
assign	pout13 = pin5;
assign	pout14 = pin18;
assign	pout15 = pin31;
assign	pout16 = pin10;
assign	pout17 = pin2;
assign	pout18 = pin8;
assign	pout19 = pin24;
assign	pout20 = pin14;
assign	pout21 = pin32;
assign	pout22 = pin27;
assign	pout23 = pin3;
assign	pout24 = pin9;
assign	pout25 = pin19;
assign	pout26 = pin13;
assign	pout27 = pin30;
assign	pout28 = pin6;
assign	pout29 = pin22;
assign	pout30 = pin11;
assign	pout31 = pin4;
assign	pout32 = pin25;




endmodule
