// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Thu Nov 25 22:52:34 2021"

module desencrypt(
	clk,
	rst_n,
	initial_key,
	reg13,
	reg12,
	reg11,
	reg10,
	reg103,
	reg102,
	reg101,
	reg100,
	reg113,
	reg112,
	reg111,
	reg110,
	reg123,
	reg122,
	reg121,
	reg120,
	reg133,
	reg132,
	reg131,
	reg130,
	reg14,
	reg15,
	reg16,
	reg2,
	reg3,
	reg4,
	reg5,
	reg6,
	reg7,
	reg8,
	reg9,
	des_encrypt_out
);


input wire	clk;
input wire	rst_n;
input wire	[63:0] initial_key;
input wire	reg13;
input wire	reg12;
input wire	reg11;
input wire	reg10;
input wire	reg103;
input wire	reg102;
input wire	reg101;
input wire	reg100;
input wire	reg113;
input wire	reg112;
input wire	reg111;
input wire	reg110;
input wire	reg123;
input wire	reg122;
input wire	reg121;
input wire	reg120;
input wire	reg133;
input wire	reg132;
input wire	reg131;
input wire	reg130;
input wire	[3:0] reg14;
input wire	[3:0] reg15;
input wire	[3:0] reg16;
input wire	[3:0] reg2;
input wire	[3:0] reg3;
input wire	[3:0] reg4;
input wire	[3:0] reg5;
input wire	[3:0] reg6;
input wire	[3:0] reg7;
input wire	[3:0] reg8;
input wire	[3:0] reg9;
output wire	[63:0] des_encrypt_out;

wire	[63:0] des_encrypt_out_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	[47:0] SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_116;
wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_128;
wire	[47:0] SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_148;
wire	SYNTHESIZED_WIRE_149;
wire	SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_151;
wire	SYNTHESIZED_WIRE_152;
wire	SYNTHESIZED_WIRE_153;
wire	SYNTHESIZED_WIRE_154;
wire	SYNTHESIZED_WIRE_155;
wire	SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_157;
wire	SYNTHESIZED_WIRE_158;
wire	SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_161;
wire	SYNTHESIZED_WIRE_162;
wire	SYNTHESIZED_WIRE_163;
wire	SYNTHESIZED_WIRE_164;
wire	SYNTHESIZED_WIRE_165;
wire	SYNTHESIZED_WIRE_166;
wire	SYNTHESIZED_WIRE_167;
wire	SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_170;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	SYNTHESIZED_WIRE_173;
wire	SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_175;
wire	SYNTHESIZED_WIRE_176;
wire	SYNTHESIZED_WIRE_177;
wire	SYNTHESIZED_WIRE_178;
wire	SYNTHESIZED_WIRE_179;
wire	SYNTHESIZED_WIRE_180;
wire	SYNTHESIZED_WIRE_181;
wire	SYNTHESIZED_WIRE_182;
wire	SYNTHESIZED_WIRE_183;
wire	SYNTHESIZED_WIRE_184;
wire	SYNTHESIZED_WIRE_185;
wire	SYNTHESIZED_WIRE_186;
wire	SYNTHESIZED_WIRE_187;
wire	SYNTHESIZED_WIRE_188;
wire	SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	SYNTHESIZED_WIRE_191;
wire	SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_193;
wire	[47:0] SYNTHESIZED_WIRE_194;
wire	SYNTHESIZED_WIRE_195;
wire	SYNTHESIZED_WIRE_196;
wire	SYNTHESIZED_WIRE_197;
wire	SYNTHESIZED_WIRE_198;
wire	SYNTHESIZED_WIRE_199;
wire	SYNTHESIZED_WIRE_200;
wire	SYNTHESIZED_WIRE_201;
wire	SYNTHESIZED_WIRE_202;
wire	SYNTHESIZED_WIRE_203;
wire	SYNTHESIZED_WIRE_204;
wire	SYNTHESIZED_WIRE_205;
wire	SYNTHESIZED_WIRE_206;
wire	SYNTHESIZED_WIRE_207;
wire	SYNTHESIZED_WIRE_208;
wire	SYNTHESIZED_WIRE_209;
wire	SYNTHESIZED_WIRE_210;
wire	SYNTHESIZED_WIRE_211;
wire	SYNTHESIZED_WIRE_212;
wire	SYNTHESIZED_WIRE_213;
wire	SYNTHESIZED_WIRE_214;
wire	SYNTHESIZED_WIRE_215;
wire	SYNTHESIZED_WIRE_216;
wire	SYNTHESIZED_WIRE_217;
wire	SYNTHESIZED_WIRE_218;
wire	SYNTHESIZED_WIRE_219;
wire	SYNTHESIZED_WIRE_220;
wire	SYNTHESIZED_WIRE_221;
wire	SYNTHESIZED_WIRE_222;
wire	SYNTHESIZED_WIRE_223;
wire	SYNTHESIZED_WIRE_224;
wire	SYNTHESIZED_WIRE_225;
wire	SYNTHESIZED_WIRE_226;
wire	SYNTHESIZED_WIRE_227;
wire	SYNTHESIZED_WIRE_228;
wire	SYNTHESIZED_WIRE_229;
wire	SYNTHESIZED_WIRE_230;
wire	SYNTHESIZED_WIRE_231;
wire	SYNTHESIZED_WIRE_232;
wire	SYNTHESIZED_WIRE_233;
wire	SYNTHESIZED_WIRE_234;
wire	SYNTHESIZED_WIRE_235;
wire	SYNTHESIZED_WIRE_236;
wire	SYNTHESIZED_WIRE_237;
wire	SYNTHESIZED_WIRE_238;
wire	SYNTHESIZED_WIRE_239;
wire	SYNTHESIZED_WIRE_240;
wire	SYNTHESIZED_WIRE_241;
wire	SYNTHESIZED_WIRE_242;
wire	SYNTHESIZED_WIRE_243;
wire	SYNTHESIZED_WIRE_244;
wire	SYNTHESIZED_WIRE_245;
wire	SYNTHESIZED_WIRE_246;
wire	SYNTHESIZED_WIRE_247;
wire	SYNTHESIZED_WIRE_248;
wire	SYNTHESIZED_WIRE_249;
wire	SYNTHESIZED_WIRE_250;
wire	SYNTHESIZED_WIRE_251;
wire	SYNTHESIZED_WIRE_252;
wire	SYNTHESIZED_WIRE_253;
wire	SYNTHESIZED_WIRE_254;
wire	SYNTHESIZED_WIRE_255;
wire	SYNTHESIZED_WIRE_256;
wire	SYNTHESIZED_WIRE_257;
wire	SYNTHESIZED_WIRE_258;
wire	SYNTHESIZED_WIRE_259;
wire	SYNTHESIZED_WIRE_260;
wire	SYNTHESIZED_WIRE_261;
wire	SYNTHESIZED_WIRE_262;
wire	SYNTHESIZED_WIRE_263;
wire	SYNTHESIZED_WIRE_264;
wire	SYNTHESIZED_WIRE_265;
wire	SYNTHESIZED_WIRE_266;
wire	SYNTHESIZED_WIRE_267;
wire	SYNTHESIZED_WIRE_268;
wire	SYNTHESIZED_WIRE_269;
wire	SYNTHESIZED_WIRE_270;
wire	SYNTHESIZED_WIRE_271;
wire	SYNTHESIZED_WIRE_272;
wire	SYNTHESIZED_WIRE_273;
wire	SYNTHESIZED_WIRE_274;
wire	SYNTHESIZED_WIRE_275;
wire	SYNTHESIZED_WIRE_276;
wire	SYNTHESIZED_WIRE_277;
wire	SYNTHESIZED_WIRE_278;
wire	SYNTHESIZED_WIRE_279;
wire	SYNTHESIZED_WIRE_280;
wire	SYNTHESIZED_WIRE_281;
wire	SYNTHESIZED_WIRE_282;
wire	SYNTHESIZED_WIRE_283;
wire	SYNTHESIZED_WIRE_284;
wire	SYNTHESIZED_WIRE_285;
wire	SYNTHESIZED_WIRE_286;
wire	SYNTHESIZED_WIRE_287;
wire	SYNTHESIZED_WIRE_288;
wire	SYNTHESIZED_WIRE_289;
wire	SYNTHESIZED_WIRE_290;
wire	SYNTHESIZED_WIRE_291;
wire	SYNTHESIZED_WIRE_292;
wire	SYNTHESIZED_WIRE_293;
wire	SYNTHESIZED_WIRE_294;
wire	SYNTHESIZED_WIRE_295;
wire	SYNTHESIZED_WIRE_296;
wire	SYNTHESIZED_WIRE_297;
wire	SYNTHESIZED_WIRE_298;
wire	SYNTHESIZED_WIRE_299;
wire	SYNTHESIZED_WIRE_300;
wire	SYNTHESIZED_WIRE_301;
wire	SYNTHESIZED_WIRE_302;
wire	SYNTHESIZED_WIRE_303;
wire	SYNTHESIZED_WIRE_304;
wire	SYNTHESIZED_WIRE_305;
wire	SYNTHESIZED_WIRE_306;
wire	SYNTHESIZED_WIRE_307;
wire	SYNTHESIZED_WIRE_308;
wire	SYNTHESIZED_WIRE_309;
wire	SYNTHESIZED_WIRE_310;
wire	SYNTHESIZED_WIRE_311;
wire	SYNTHESIZED_WIRE_312;
wire	SYNTHESIZED_WIRE_313;
wire	SYNTHESIZED_WIRE_314;
wire	SYNTHESIZED_WIRE_315;
wire	SYNTHESIZED_WIRE_316;
wire	SYNTHESIZED_WIRE_317;
wire	SYNTHESIZED_WIRE_318;
wire	SYNTHESIZED_WIRE_319;
wire	SYNTHESIZED_WIRE_320;
wire	SYNTHESIZED_WIRE_321;
wire	SYNTHESIZED_WIRE_322;
wire	[47:0] SYNTHESIZED_WIRE_323;
wire	SYNTHESIZED_WIRE_324;
wire	SYNTHESIZED_WIRE_325;
wire	SYNTHESIZED_WIRE_326;
wire	SYNTHESIZED_WIRE_327;
wire	SYNTHESIZED_WIRE_328;
wire	SYNTHESIZED_WIRE_329;
wire	SYNTHESIZED_WIRE_330;
wire	SYNTHESIZED_WIRE_331;
wire	SYNTHESIZED_WIRE_332;
wire	SYNTHESIZED_WIRE_333;
wire	SYNTHESIZED_WIRE_334;
wire	SYNTHESIZED_WIRE_335;
wire	SYNTHESIZED_WIRE_336;
wire	SYNTHESIZED_WIRE_337;
wire	SYNTHESIZED_WIRE_338;
wire	SYNTHESIZED_WIRE_339;
wire	SYNTHESIZED_WIRE_340;
wire	SYNTHESIZED_WIRE_341;
wire	SYNTHESIZED_WIRE_342;
wire	SYNTHESIZED_WIRE_343;
wire	SYNTHESIZED_WIRE_344;
wire	SYNTHESIZED_WIRE_345;
wire	SYNTHESIZED_WIRE_346;
wire	SYNTHESIZED_WIRE_347;
wire	SYNTHESIZED_WIRE_348;
wire	SYNTHESIZED_WIRE_349;
wire	SYNTHESIZED_WIRE_350;
wire	SYNTHESIZED_WIRE_351;
wire	SYNTHESIZED_WIRE_352;
wire	SYNTHESIZED_WIRE_353;
wire	SYNTHESIZED_WIRE_354;
wire	SYNTHESIZED_WIRE_355;
wire	SYNTHESIZED_WIRE_356;
wire	SYNTHESIZED_WIRE_357;
wire	SYNTHESIZED_WIRE_358;
wire	SYNTHESIZED_WIRE_359;
wire	SYNTHESIZED_WIRE_360;
wire	SYNTHESIZED_WIRE_361;
wire	SYNTHESIZED_WIRE_362;
wire	SYNTHESIZED_WIRE_363;
wire	SYNTHESIZED_WIRE_364;
wire	SYNTHESIZED_WIRE_365;
wire	SYNTHESIZED_WIRE_366;
wire	SYNTHESIZED_WIRE_367;
wire	SYNTHESIZED_WIRE_368;
wire	SYNTHESIZED_WIRE_369;
wire	SYNTHESIZED_WIRE_370;
wire	SYNTHESIZED_WIRE_371;
wire	SYNTHESIZED_WIRE_372;
wire	SYNTHESIZED_WIRE_373;
wire	SYNTHESIZED_WIRE_374;
wire	SYNTHESIZED_WIRE_375;
wire	SYNTHESIZED_WIRE_376;
wire	SYNTHESIZED_WIRE_377;
wire	SYNTHESIZED_WIRE_378;
wire	SYNTHESIZED_WIRE_379;
wire	SYNTHESIZED_WIRE_380;
wire	SYNTHESIZED_WIRE_381;
wire	SYNTHESIZED_WIRE_382;
wire	SYNTHESIZED_WIRE_383;
wire	SYNTHESIZED_WIRE_384;
wire	SYNTHESIZED_WIRE_385;
wire	SYNTHESIZED_WIRE_386;
wire	SYNTHESIZED_WIRE_387;
wire	[47:0] SYNTHESIZED_WIRE_388;
wire	SYNTHESIZED_WIRE_389;
wire	SYNTHESIZED_WIRE_390;
wire	SYNTHESIZED_WIRE_391;
wire	SYNTHESIZED_WIRE_392;
wire	SYNTHESIZED_WIRE_393;
wire	SYNTHESIZED_WIRE_394;
wire	SYNTHESIZED_WIRE_395;
wire	SYNTHESIZED_WIRE_396;
wire	SYNTHESIZED_WIRE_397;
wire	SYNTHESIZED_WIRE_398;
wire	SYNTHESIZED_WIRE_399;
wire	SYNTHESIZED_WIRE_400;
wire	SYNTHESIZED_WIRE_401;
wire	SYNTHESIZED_WIRE_402;
wire	SYNTHESIZED_WIRE_403;
wire	SYNTHESIZED_WIRE_404;
wire	SYNTHESIZED_WIRE_405;
wire	SYNTHESIZED_WIRE_406;
wire	SYNTHESIZED_WIRE_407;
wire	SYNTHESIZED_WIRE_408;
wire	SYNTHESIZED_WIRE_409;
wire	SYNTHESIZED_WIRE_410;
wire	SYNTHESIZED_WIRE_411;
wire	SYNTHESIZED_WIRE_412;
wire	SYNTHESIZED_WIRE_413;
wire	SYNTHESIZED_WIRE_414;
wire	SYNTHESIZED_WIRE_415;
wire	SYNTHESIZED_WIRE_416;
wire	SYNTHESIZED_WIRE_417;
wire	SYNTHESIZED_WIRE_418;
wire	SYNTHESIZED_WIRE_419;
wire	SYNTHESIZED_WIRE_420;
wire	SYNTHESIZED_WIRE_421;
wire	SYNTHESIZED_WIRE_422;
wire	SYNTHESIZED_WIRE_423;
wire	SYNTHESIZED_WIRE_424;
wire	SYNTHESIZED_WIRE_425;
wire	SYNTHESIZED_WIRE_426;
wire	SYNTHESIZED_WIRE_427;
wire	SYNTHESIZED_WIRE_428;
wire	SYNTHESIZED_WIRE_429;
wire	SYNTHESIZED_WIRE_430;
wire	SYNTHESIZED_WIRE_431;
wire	SYNTHESIZED_WIRE_432;
wire	SYNTHESIZED_WIRE_433;
wire	SYNTHESIZED_WIRE_434;
wire	SYNTHESIZED_WIRE_435;
wire	SYNTHESIZED_WIRE_436;
wire	SYNTHESIZED_WIRE_437;
wire	SYNTHESIZED_WIRE_438;
wire	SYNTHESIZED_WIRE_439;
wire	SYNTHESIZED_WIRE_440;
wire	SYNTHESIZED_WIRE_441;
wire	SYNTHESIZED_WIRE_442;
wire	SYNTHESIZED_WIRE_443;
wire	SYNTHESIZED_WIRE_444;
wire	SYNTHESIZED_WIRE_445;
wire	SYNTHESIZED_WIRE_446;
wire	SYNTHESIZED_WIRE_447;
wire	SYNTHESIZED_WIRE_448;
wire	SYNTHESIZED_WIRE_449;
wire	SYNTHESIZED_WIRE_450;
wire	SYNTHESIZED_WIRE_451;
wire	SYNTHESIZED_WIRE_452;
wire	[47:0] SYNTHESIZED_WIRE_453;
wire	SYNTHESIZED_WIRE_454;
wire	SYNTHESIZED_WIRE_455;
wire	SYNTHESIZED_WIRE_456;
wire	SYNTHESIZED_WIRE_457;
wire	SYNTHESIZED_WIRE_458;
wire	SYNTHESIZED_WIRE_459;
wire	SYNTHESIZED_WIRE_460;
wire	SYNTHESIZED_WIRE_461;
wire	SYNTHESIZED_WIRE_462;
wire	SYNTHESIZED_WIRE_463;
wire	SYNTHESIZED_WIRE_464;
wire	SYNTHESIZED_WIRE_465;
wire	SYNTHESIZED_WIRE_466;
wire	SYNTHESIZED_WIRE_467;
wire	SYNTHESIZED_WIRE_468;
wire	SYNTHESIZED_WIRE_469;
wire	SYNTHESIZED_WIRE_470;
wire	SYNTHESIZED_WIRE_471;
wire	SYNTHESIZED_WIRE_472;
wire	SYNTHESIZED_WIRE_473;
wire	SYNTHESIZED_WIRE_474;
wire	SYNTHESIZED_WIRE_475;
wire	SYNTHESIZED_WIRE_476;
wire	SYNTHESIZED_WIRE_477;
wire	SYNTHESIZED_WIRE_478;
wire	SYNTHESIZED_WIRE_479;
wire	SYNTHESIZED_WIRE_480;
wire	SYNTHESIZED_WIRE_481;
wire	SYNTHESIZED_WIRE_482;
wire	SYNTHESIZED_WIRE_483;
wire	SYNTHESIZED_WIRE_484;
wire	SYNTHESIZED_WIRE_485;
wire	SYNTHESIZED_WIRE_486;
wire	SYNTHESIZED_WIRE_487;
wire	SYNTHESIZED_WIRE_488;
wire	SYNTHESIZED_WIRE_489;
wire	SYNTHESIZED_WIRE_490;
wire	SYNTHESIZED_WIRE_491;
wire	SYNTHESIZED_WIRE_492;
wire	SYNTHESIZED_WIRE_493;
wire	SYNTHESIZED_WIRE_494;
wire	SYNTHESIZED_WIRE_495;
wire	SYNTHESIZED_WIRE_496;
wire	SYNTHESIZED_WIRE_497;
wire	SYNTHESIZED_WIRE_498;
wire	SYNTHESIZED_WIRE_499;
wire	SYNTHESIZED_WIRE_500;
wire	SYNTHESIZED_WIRE_501;
wire	SYNTHESIZED_WIRE_502;
wire	SYNTHESIZED_WIRE_503;
wire	SYNTHESIZED_WIRE_504;
wire	SYNTHESIZED_WIRE_505;
wire	SYNTHESIZED_WIRE_506;
wire	SYNTHESIZED_WIRE_507;
wire	SYNTHESIZED_WIRE_508;
wire	SYNTHESIZED_WIRE_509;
wire	SYNTHESIZED_WIRE_510;
wire	SYNTHESIZED_WIRE_511;
wire	SYNTHESIZED_WIRE_512;
wire	SYNTHESIZED_WIRE_513;
wire	SYNTHESIZED_WIRE_514;
wire	SYNTHESIZED_WIRE_515;
wire	SYNTHESIZED_WIRE_516;
wire	SYNTHESIZED_WIRE_517;
wire	[47:0] SYNTHESIZED_WIRE_518;
wire	SYNTHESIZED_WIRE_519;
wire	SYNTHESIZED_WIRE_520;
wire	SYNTHESIZED_WIRE_521;
wire	SYNTHESIZED_WIRE_522;
wire	SYNTHESIZED_WIRE_523;
wire	SYNTHESIZED_WIRE_524;
wire	SYNTHESIZED_WIRE_525;
wire	SYNTHESIZED_WIRE_526;
wire	SYNTHESIZED_WIRE_527;
wire	SYNTHESIZED_WIRE_528;
wire	SYNTHESIZED_WIRE_529;
wire	SYNTHESIZED_WIRE_530;
wire	SYNTHESIZED_WIRE_531;
wire	SYNTHESIZED_WIRE_532;
wire	SYNTHESIZED_WIRE_533;
wire	SYNTHESIZED_WIRE_534;
wire	SYNTHESIZED_WIRE_535;
wire	SYNTHESIZED_WIRE_536;
wire	SYNTHESIZED_WIRE_537;
wire	SYNTHESIZED_WIRE_538;
wire	SYNTHESIZED_WIRE_539;
wire	SYNTHESIZED_WIRE_540;
wire	SYNTHESIZED_WIRE_541;
wire	SYNTHESIZED_WIRE_542;
wire	SYNTHESIZED_WIRE_543;
wire	SYNTHESIZED_WIRE_544;
wire	SYNTHESIZED_WIRE_545;
wire	SYNTHESIZED_WIRE_546;
wire	SYNTHESIZED_WIRE_547;
wire	SYNTHESIZED_WIRE_548;
wire	SYNTHESIZED_WIRE_549;
wire	SYNTHESIZED_WIRE_550;
wire	SYNTHESIZED_WIRE_551;
wire	SYNTHESIZED_WIRE_552;
wire	SYNTHESIZED_WIRE_553;
wire	SYNTHESIZED_WIRE_554;
wire	SYNTHESIZED_WIRE_555;
wire	SYNTHESIZED_WIRE_556;
wire	SYNTHESIZED_WIRE_557;
wire	SYNTHESIZED_WIRE_558;
wire	SYNTHESIZED_WIRE_559;
wire	SYNTHESIZED_WIRE_560;
wire	SYNTHESIZED_WIRE_561;
wire	SYNTHESIZED_WIRE_562;
wire	SYNTHESIZED_WIRE_563;
wire	SYNTHESIZED_WIRE_564;
wire	SYNTHESIZED_WIRE_565;
wire	SYNTHESIZED_WIRE_566;
wire	SYNTHESIZED_WIRE_567;
wire	SYNTHESIZED_WIRE_568;
wire	SYNTHESIZED_WIRE_569;
wire	SYNTHESIZED_WIRE_570;
wire	SYNTHESIZED_WIRE_571;
wire	SYNTHESIZED_WIRE_572;
wire	SYNTHESIZED_WIRE_573;
wire	SYNTHESIZED_WIRE_574;
wire	SYNTHESIZED_WIRE_575;
wire	SYNTHESIZED_WIRE_576;
wire	SYNTHESIZED_WIRE_577;
wire	SYNTHESIZED_WIRE_578;
wire	SYNTHESIZED_WIRE_579;
wire	SYNTHESIZED_WIRE_580;
wire	SYNTHESIZED_WIRE_581;
wire	SYNTHESIZED_WIRE_582;
wire	[47:0] SYNTHESIZED_WIRE_583;
wire	SYNTHESIZED_WIRE_584;
wire	SYNTHESIZED_WIRE_585;
wire	SYNTHESIZED_WIRE_586;
wire	SYNTHESIZED_WIRE_587;
wire	SYNTHESIZED_WIRE_588;
wire	SYNTHESIZED_WIRE_589;
wire	SYNTHESIZED_WIRE_590;
wire	SYNTHESIZED_WIRE_591;
wire	SYNTHESIZED_WIRE_592;
wire	SYNTHESIZED_WIRE_593;
wire	SYNTHESIZED_WIRE_594;
wire	SYNTHESIZED_WIRE_595;
wire	SYNTHESIZED_WIRE_596;
wire	SYNTHESIZED_WIRE_597;
wire	SYNTHESIZED_WIRE_598;
wire	SYNTHESIZED_WIRE_599;
wire	SYNTHESIZED_WIRE_600;
wire	SYNTHESIZED_WIRE_601;
wire	SYNTHESIZED_WIRE_602;
wire	SYNTHESIZED_WIRE_603;
wire	SYNTHESIZED_WIRE_604;
wire	SYNTHESIZED_WIRE_605;
wire	SYNTHESIZED_WIRE_606;
wire	SYNTHESIZED_WIRE_607;
wire	SYNTHESIZED_WIRE_608;
wire	SYNTHESIZED_WIRE_609;
wire	SYNTHESIZED_WIRE_610;
wire	SYNTHESIZED_WIRE_611;
wire	SYNTHESIZED_WIRE_612;
wire	SYNTHESIZED_WIRE_613;
wire	SYNTHESIZED_WIRE_614;
wire	SYNTHESIZED_WIRE_615;
wire	SYNTHESIZED_WIRE_616;
wire	SYNTHESIZED_WIRE_617;
wire	SYNTHESIZED_WIRE_618;
wire	SYNTHESIZED_WIRE_619;
wire	SYNTHESIZED_WIRE_620;
wire	SYNTHESIZED_WIRE_621;
wire	SYNTHESIZED_WIRE_622;
wire	SYNTHESIZED_WIRE_623;
wire	SYNTHESIZED_WIRE_624;
wire	SYNTHESIZED_WIRE_625;
wire	SYNTHESIZED_WIRE_626;
wire	SYNTHESIZED_WIRE_627;
wire	SYNTHESIZED_WIRE_628;
wire	SYNTHESIZED_WIRE_629;
wire	SYNTHESIZED_WIRE_630;
wire	SYNTHESIZED_WIRE_631;
wire	SYNTHESIZED_WIRE_632;
wire	SYNTHESIZED_WIRE_633;
wire	SYNTHESIZED_WIRE_634;
wire	SYNTHESIZED_WIRE_635;
wire	SYNTHESIZED_WIRE_636;
wire	SYNTHESIZED_WIRE_637;
wire	SYNTHESIZED_WIRE_638;
wire	SYNTHESIZED_WIRE_639;
wire	SYNTHESIZED_WIRE_640;
wire	SYNTHESIZED_WIRE_641;
wire	SYNTHESIZED_WIRE_642;
wire	SYNTHESIZED_WIRE_643;
wire	SYNTHESIZED_WIRE_644;
wire	SYNTHESIZED_WIRE_645;
wire	SYNTHESIZED_WIRE_646;
wire	SYNTHESIZED_WIRE_647;
wire	[47:0] SYNTHESIZED_WIRE_648;
wire	SYNTHESIZED_WIRE_649;
wire	SYNTHESIZED_WIRE_650;
wire	SYNTHESIZED_WIRE_651;
wire	SYNTHESIZED_WIRE_652;
wire	SYNTHESIZED_WIRE_653;
wire	SYNTHESIZED_WIRE_654;
wire	SYNTHESIZED_WIRE_655;
wire	SYNTHESIZED_WIRE_656;
wire	SYNTHESIZED_WIRE_657;
wire	SYNTHESIZED_WIRE_658;
wire	SYNTHESIZED_WIRE_659;
wire	SYNTHESIZED_WIRE_660;
wire	SYNTHESIZED_WIRE_661;
wire	SYNTHESIZED_WIRE_662;
wire	SYNTHESIZED_WIRE_663;
wire	SYNTHESIZED_WIRE_664;
wire	SYNTHESIZED_WIRE_665;
wire	SYNTHESIZED_WIRE_666;
wire	SYNTHESIZED_WIRE_667;
wire	SYNTHESIZED_WIRE_668;
wire	SYNTHESIZED_WIRE_669;
wire	SYNTHESIZED_WIRE_670;
wire	SYNTHESIZED_WIRE_671;
wire	SYNTHESIZED_WIRE_672;
wire	SYNTHESIZED_WIRE_673;
wire	SYNTHESIZED_WIRE_674;
wire	SYNTHESIZED_WIRE_675;
wire	SYNTHESIZED_WIRE_676;
wire	SYNTHESIZED_WIRE_677;
wire	SYNTHESIZED_WIRE_678;
wire	SYNTHESIZED_WIRE_679;
wire	SYNTHESIZED_WIRE_680;
wire	SYNTHESIZED_WIRE_681;
wire	SYNTHESIZED_WIRE_682;
wire	SYNTHESIZED_WIRE_683;
wire	SYNTHESIZED_WIRE_684;
wire	SYNTHESIZED_WIRE_685;
wire	SYNTHESIZED_WIRE_686;
wire	SYNTHESIZED_WIRE_687;
wire	SYNTHESIZED_WIRE_688;
wire	SYNTHESIZED_WIRE_689;
wire	SYNTHESIZED_WIRE_690;
wire	SYNTHESIZED_WIRE_691;
wire	SYNTHESIZED_WIRE_692;
wire	SYNTHESIZED_WIRE_693;
wire	SYNTHESIZED_WIRE_694;
wire	SYNTHESIZED_WIRE_695;
wire	SYNTHESIZED_WIRE_696;
wire	SYNTHESIZED_WIRE_697;
wire	SYNTHESIZED_WIRE_698;
wire	SYNTHESIZED_WIRE_699;
wire	SYNTHESIZED_WIRE_700;
wire	SYNTHESIZED_WIRE_701;
wire	SYNTHESIZED_WIRE_702;
wire	SYNTHESIZED_WIRE_703;
wire	SYNTHESIZED_WIRE_704;
wire	SYNTHESIZED_WIRE_705;
wire	SYNTHESIZED_WIRE_706;
wire	SYNTHESIZED_WIRE_707;
wire	SYNTHESIZED_WIRE_708;
wire	SYNTHESIZED_WIRE_709;
wire	SYNTHESIZED_WIRE_710;
wire	SYNTHESIZED_WIRE_711;
wire	SYNTHESIZED_WIRE_712;
wire	[47:0] SYNTHESIZED_WIRE_713;
wire	SYNTHESIZED_WIRE_714;
wire	SYNTHESIZED_WIRE_715;
wire	SYNTHESIZED_WIRE_716;
wire	SYNTHESIZED_WIRE_717;
wire	SYNTHESIZED_WIRE_718;
wire	SYNTHESIZED_WIRE_719;
wire	SYNTHESIZED_WIRE_720;
wire	SYNTHESIZED_WIRE_721;
wire	SYNTHESIZED_WIRE_722;
wire	SYNTHESIZED_WIRE_723;
wire	SYNTHESIZED_WIRE_724;
wire	SYNTHESIZED_WIRE_725;
wire	SYNTHESIZED_WIRE_726;
wire	SYNTHESIZED_WIRE_727;
wire	SYNTHESIZED_WIRE_728;
wire	SYNTHESIZED_WIRE_729;
wire	SYNTHESIZED_WIRE_730;
wire	SYNTHESIZED_WIRE_731;
wire	SYNTHESIZED_WIRE_732;
wire	SYNTHESIZED_WIRE_733;
wire	SYNTHESIZED_WIRE_734;
wire	SYNTHESIZED_WIRE_735;
wire	SYNTHESIZED_WIRE_736;
wire	SYNTHESIZED_WIRE_737;
wire	SYNTHESIZED_WIRE_738;
wire	SYNTHESIZED_WIRE_739;
wire	SYNTHESIZED_WIRE_740;
wire	SYNTHESIZED_WIRE_741;
wire	SYNTHESIZED_WIRE_742;
wire	SYNTHESIZED_WIRE_743;
wire	SYNTHESIZED_WIRE_744;
wire	SYNTHESIZED_WIRE_745;
wire	SYNTHESIZED_WIRE_746;
wire	SYNTHESIZED_WIRE_747;
wire	SYNTHESIZED_WIRE_748;
wire	SYNTHESIZED_WIRE_749;
wire	SYNTHESIZED_WIRE_750;
wire	SYNTHESIZED_WIRE_751;
wire	SYNTHESIZED_WIRE_752;
wire	SYNTHESIZED_WIRE_753;
wire	SYNTHESIZED_WIRE_754;
wire	SYNTHESIZED_WIRE_755;
wire	SYNTHESIZED_WIRE_756;
wire	SYNTHESIZED_WIRE_757;
wire	SYNTHESIZED_WIRE_758;
wire	SYNTHESIZED_WIRE_759;
wire	SYNTHESIZED_WIRE_760;
wire	SYNTHESIZED_WIRE_761;
wire	SYNTHESIZED_WIRE_762;
wire	SYNTHESIZED_WIRE_763;
wire	SYNTHESIZED_WIRE_764;
wire	SYNTHESIZED_WIRE_765;
wire	SYNTHESIZED_WIRE_766;
wire	SYNTHESIZED_WIRE_767;
wire	SYNTHESIZED_WIRE_768;
wire	SYNTHESIZED_WIRE_769;
wire	SYNTHESIZED_WIRE_770;
wire	SYNTHESIZED_WIRE_771;
wire	SYNTHESIZED_WIRE_772;
wire	SYNTHESIZED_WIRE_773;
wire	SYNTHESIZED_WIRE_774;
wire	SYNTHESIZED_WIRE_775;
wire	SYNTHESIZED_WIRE_776;
wire	SYNTHESIZED_WIRE_777;
wire	[47:0] SYNTHESIZED_WIRE_778;
wire	SYNTHESIZED_WIRE_779;
wire	SYNTHESIZED_WIRE_780;
wire	SYNTHESIZED_WIRE_781;
wire	SYNTHESIZED_WIRE_782;
wire	SYNTHESIZED_WIRE_783;
wire	SYNTHESIZED_WIRE_784;
wire	SYNTHESIZED_WIRE_785;
wire	SYNTHESIZED_WIRE_786;
wire	SYNTHESIZED_WIRE_787;
wire	SYNTHESIZED_WIRE_788;
wire	SYNTHESIZED_WIRE_789;
wire	SYNTHESIZED_WIRE_790;
wire	SYNTHESIZED_WIRE_791;
wire	SYNTHESIZED_WIRE_792;
wire	SYNTHESIZED_WIRE_793;
wire	SYNTHESIZED_WIRE_794;
wire	SYNTHESIZED_WIRE_795;
wire	SYNTHESIZED_WIRE_796;
wire	SYNTHESIZED_WIRE_797;
wire	SYNTHESIZED_WIRE_798;
wire	SYNTHESIZED_WIRE_799;
wire	SYNTHESIZED_WIRE_800;
wire	SYNTHESIZED_WIRE_801;
wire	SYNTHESIZED_WIRE_802;
wire	SYNTHESIZED_WIRE_803;
wire	SYNTHESIZED_WIRE_804;
wire	SYNTHESIZED_WIRE_805;
wire	SYNTHESIZED_WIRE_806;
wire	SYNTHESIZED_WIRE_807;
wire	SYNTHESIZED_WIRE_808;
wire	SYNTHESIZED_WIRE_809;
wire	SYNTHESIZED_WIRE_810;
wire	SYNTHESIZED_WIRE_811;
wire	SYNTHESIZED_WIRE_812;
wire	SYNTHESIZED_WIRE_813;
wire	SYNTHESIZED_WIRE_814;
wire	SYNTHESIZED_WIRE_815;
wire	SYNTHESIZED_WIRE_816;
wire	SYNTHESIZED_WIRE_817;
wire	SYNTHESIZED_WIRE_818;
wire	SYNTHESIZED_WIRE_819;
wire	SYNTHESIZED_WIRE_820;
wire	SYNTHESIZED_WIRE_821;
wire	SYNTHESIZED_WIRE_822;
wire	SYNTHESIZED_WIRE_823;
wire	SYNTHESIZED_WIRE_824;
wire	SYNTHESIZED_WIRE_825;
wire	SYNTHESIZED_WIRE_826;
wire	SYNTHESIZED_WIRE_827;
wire	SYNTHESIZED_WIRE_828;
wire	SYNTHESIZED_WIRE_829;
wire	SYNTHESIZED_WIRE_830;
wire	SYNTHESIZED_WIRE_831;
wire	SYNTHESIZED_WIRE_832;
wire	SYNTHESIZED_WIRE_833;
wire	SYNTHESIZED_WIRE_834;
wire	SYNTHESIZED_WIRE_835;
wire	SYNTHESIZED_WIRE_836;
wire	SYNTHESIZED_WIRE_837;
wire	SYNTHESIZED_WIRE_838;
wire	SYNTHESIZED_WIRE_839;
wire	SYNTHESIZED_WIRE_840;
wire	SYNTHESIZED_WIRE_841;
wire	SYNTHESIZED_WIRE_842;
wire	[47:0] SYNTHESIZED_WIRE_843;
wire	SYNTHESIZED_WIRE_844;
wire	SYNTHESIZED_WIRE_845;
wire	SYNTHESIZED_WIRE_846;
wire	SYNTHESIZED_WIRE_847;
wire	SYNTHESIZED_WIRE_848;
wire	SYNTHESIZED_WIRE_849;
wire	SYNTHESIZED_WIRE_850;
wire	SYNTHESIZED_WIRE_851;
wire	SYNTHESIZED_WIRE_852;
wire	SYNTHESIZED_WIRE_853;
wire	SYNTHESIZED_WIRE_854;
wire	SYNTHESIZED_WIRE_855;
wire	SYNTHESIZED_WIRE_856;
wire	SYNTHESIZED_WIRE_857;
wire	SYNTHESIZED_WIRE_858;
wire	SYNTHESIZED_WIRE_859;
wire	SYNTHESIZED_WIRE_860;
wire	SYNTHESIZED_WIRE_861;
wire	SYNTHESIZED_WIRE_862;
wire	SYNTHESIZED_WIRE_863;
wire	SYNTHESIZED_WIRE_864;
wire	SYNTHESIZED_WIRE_865;
wire	SYNTHESIZED_WIRE_866;
wire	SYNTHESIZED_WIRE_867;
wire	SYNTHESIZED_WIRE_868;
wire	SYNTHESIZED_WIRE_869;
wire	SYNTHESIZED_WIRE_870;
wire	SYNTHESIZED_WIRE_871;
wire	SYNTHESIZED_WIRE_872;
wire	SYNTHESIZED_WIRE_873;
wire	SYNTHESIZED_WIRE_874;
wire	SYNTHESIZED_WIRE_875;
wire	SYNTHESIZED_WIRE_876;
wire	SYNTHESIZED_WIRE_877;
wire	SYNTHESIZED_WIRE_878;
wire	SYNTHESIZED_WIRE_879;
wire	SYNTHESIZED_WIRE_880;
wire	SYNTHESIZED_WIRE_881;
wire	SYNTHESIZED_WIRE_882;
wire	SYNTHESIZED_WIRE_883;
wire	SYNTHESIZED_WIRE_884;
wire	SYNTHESIZED_WIRE_885;
wire	SYNTHESIZED_WIRE_886;
wire	SYNTHESIZED_WIRE_887;
wire	SYNTHESIZED_WIRE_888;
wire	SYNTHESIZED_WIRE_889;
wire	SYNTHESIZED_WIRE_890;
wire	SYNTHESIZED_WIRE_891;
wire	SYNTHESIZED_WIRE_892;
wire	SYNTHESIZED_WIRE_893;
wire	SYNTHESIZED_WIRE_894;
wire	SYNTHESIZED_WIRE_895;
wire	SYNTHESIZED_WIRE_896;
wire	SYNTHESIZED_WIRE_897;
wire	SYNTHESIZED_WIRE_898;
wire	SYNTHESIZED_WIRE_899;
wire	SYNTHESIZED_WIRE_900;
wire	SYNTHESIZED_WIRE_901;
wire	SYNTHESIZED_WIRE_902;
wire	SYNTHESIZED_WIRE_903;
wire	SYNTHESIZED_WIRE_904;
wire	SYNTHESIZED_WIRE_905;
wire	SYNTHESIZED_WIRE_906;
wire	SYNTHESIZED_WIRE_907;
wire	[47:0] SYNTHESIZED_WIRE_908;
wire	SYNTHESIZED_WIRE_909;
wire	SYNTHESIZED_WIRE_910;
wire	SYNTHESIZED_WIRE_911;
wire	SYNTHESIZED_WIRE_912;
wire	SYNTHESIZED_WIRE_913;
wire	SYNTHESIZED_WIRE_914;
wire	SYNTHESIZED_WIRE_915;
wire	SYNTHESIZED_WIRE_916;
wire	SYNTHESIZED_WIRE_917;
wire	SYNTHESIZED_WIRE_918;
wire	SYNTHESIZED_WIRE_919;
wire	SYNTHESIZED_WIRE_920;
wire	SYNTHESIZED_WIRE_921;
wire	SYNTHESIZED_WIRE_922;
wire	SYNTHESIZED_WIRE_923;
wire	SYNTHESIZED_WIRE_924;
wire	SYNTHESIZED_WIRE_925;
wire	SYNTHESIZED_WIRE_926;
wire	SYNTHESIZED_WIRE_927;
wire	SYNTHESIZED_WIRE_928;
wire	SYNTHESIZED_WIRE_929;
wire	SYNTHESIZED_WIRE_930;
wire	SYNTHESIZED_WIRE_931;
wire	SYNTHESIZED_WIRE_932;
wire	SYNTHESIZED_WIRE_933;
wire	SYNTHESIZED_WIRE_934;
wire	SYNTHESIZED_WIRE_935;
wire	SYNTHESIZED_WIRE_936;
wire	SYNTHESIZED_WIRE_937;
wire	SYNTHESIZED_WIRE_938;
wire	SYNTHESIZED_WIRE_939;
wire	SYNTHESIZED_WIRE_940;
wire	SYNTHESIZED_WIRE_941;
wire	SYNTHESIZED_WIRE_942;
wire	SYNTHESIZED_WIRE_943;
wire	SYNTHESIZED_WIRE_944;
wire	SYNTHESIZED_WIRE_945;
wire	SYNTHESIZED_WIRE_946;
wire	SYNTHESIZED_WIRE_947;
wire	SYNTHESIZED_WIRE_948;
wire	SYNTHESIZED_WIRE_949;
wire	SYNTHESIZED_WIRE_950;
wire	SYNTHESIZED_WIRE_951;
wire	SYNTHESIZED_WIRE_952;
wire	SYNTHESIZED_WIRE_953;
wire	SYNTHESIZED_WIRE_954;
wire	SYNTHESIZED_WIRE_955;
wire	SYNTHESIZED_WIRE_956;
wire	SYNTHESIZED_WIRE_957;
wire	SYNTHESIZED_WIRE_958;
wire	SYNTHESIZED_WIRE_959;
wire	SYNTHESIZED_WIRE_960;
wire	SYNTHESIZED_WIRE_961;
wire	SYNTHESIZED_WIRE_962;
wire	SYNTHESIZED_WIRE_963;
wire	SYNTHESIZED_WIRE_964;
wire	SYNTHESIZED_WIRE_965;
wire	SYNTHESIZED_WIRE_966;
wire	SYNTHESIZED_WIRE_967;
wire	SYNTHESIZED_WIRE_968;
wire	SYNTHESIZED_WIRE_969;
wire	SYNTHESIZED_WIRE_970;
wire	SYNTHESIZED_WIRE_971;
wire	SYNTHESIZED_WIRE_972;
wire	[47:0] SYNTHESIZED_WIRE_973;
wire	SYNTHESIZED_WIRE_974;
wire	SYNTHESIZED_WIRE_975;
wire	SYNTHESIZED_WIRE_976;
wire	SYNTHESIZED_WIRE_977;
wire	SYNTHESIZED_WIRE_978;
wire	SYNTHESIZED_WIRE_979;
wire	SYNTHESIZED_WIRE_980;
wire	SYNTHESIZED_WIRE_981;
wire	SYNTHESIZED_WIRE_982;
wire	SYNTHESIZED_WIRE_983;
wire	SYNTHESIZED_WIRE_984;
wire	SYNTHESIZED_WIRE_985;
wire	SYNTHESIZED_WIRE_986;
wire	SYNTHESIZED_WIRE_987;
wire	SYNTHESIZED_WIRE_988;
wire	SYNTHESIZED_WIRE_989;
wire	SYNTHESIZED_WIRE_990;
wire	SYNTHESIZED_WIRE_991;
wire	SYNTHESIZED_WIRE_992;
wire	SYNTHESIZED_WIRE_993;
wire	SYNTHESIZED_WIRE_994;
wire	SYNTHESIZED_WIRE_995;
wire	SYNTHESIZED_WIRE_996;
wire	SYNTHESIZED_WIRE_997;
wire	SYNTHESIZED_WIRE_998;
wire	SYNTHESIZED_WIRE_999;
wire	SYNTHESIZED_WIRE_1000;
wire	SYNTHESIZED_WIRE_1001;
wire	SYNTHESIZED_WIRE_1002;
wire	SYNTHESIZED_WIRE_1003;
wire	SYNTHESIZED_WIRE_1004;
wire	SYNTHESIZED_WIRE_1005;
wire	SYNTHESIZED_WIRE_1006;
wire	SYNTHESIZED_WIRE_1007;
wire	SYNTHESIZED_WIRE_1008;
wire	SYNTHESIZED_WIRE_1009;
wire	SYNTHESIZED_WIRE_1010;
wire	SYNTHESIZED_WIRE_1011;
wire	SYNTHESIZED_WIRE_1012;
wire	SYNTHESIZED_WIRE_1013;
wire	SYNTHESIZED_WIRE_1014;
wire	SYNTHESIZED_WIRE_1015;
wire	SYNTHESIZED_WIRE_1016;
wire	SYNTHESIZED_WIRE_1017;
wire	SYNTHESIZED_WIRE_1018;
wire	SYNTHESIZED_WIRE_1019;
wire	SYNTHESIZED_WIRE_1020;
wire	SYNTHESIZED_WIRE_1021;
wire	SYNTHESIZED_WIRE_1022;
wire	SYNTHESIZED_WIRE_1023;
wire	SYNTHESIZED_WIRE_1024;
wire	SYNTHESIZED_WIRE_1025;
wire	SYNTHESIZED_WIRE_1026;
wire	SYNTHESIZED_WIRE_1027;
wire	SYNTHESIZED_WIRE_1028;
wire	SYNTHESIZED_WIRE_1029;
wire	SYNTHESIZED_WIRE_1030;
wire	SYNTHESIZED_WIRE_1031;
wire	SYNTHESIZED_WIRE_1032;
wire	SYNTHESIZED_WIRE_1033;
wire	SYNTHESIZED_WIRE_1034;
wire	SYNTHESIZED_WIRE_1035;
wire	SYNTHESIZED_WIRE_1036;
wire	SYNTHESIZED_WIRE_1037;
wire	[47:0] SYNTHESIZED_WIRE_1038;
wire	SYNTHESIZED_WIRE_1039;
wire	SYNTHESIZED_WIRE_1040;
wire	SYNTHESIZED_WIRE_1041;
wire	SYNTHESIZED_WIRE_1042;
wire	SYNTHESIZED_WIRE_1043;
wire	SYNTHESIZED_WIRE_1044;
wire	SYNTHESIZED_WIRE_1045;
wire	SYNTHESIZED_WIRE_1046;
wire	SYNTHESIZED_WIRE_1047;
wire	SYNTHESIZED_WIRE_1048;
wire	SYNTHESIZED_WIRE_1049;
wire	SYNTHESIZED_WIRE_1050;
wire	SYNTHESIZED_WIRE_1051;
wire	SYNTHESIZED_WIRE_1052;
wire	SYNTHESIZED_WIRE_1053;
wire	SYNTHESIZED_WIRE_1054;
wire	SYNTHESIZED_WIRE_1055;
wire	SYNTHESIZED_WIRE_1056;
wire	SYNTHESIZED_WIRE_1057;
wire	SYNTHESIZED_WIRE_1058;
wire	SYNTHESIZED_WIRE_1059;
wire	SYNTHESIZED_WIRE_1060;
wire	SYNTHESIZED_WIRE_1061;
wire	SYNTHESIZED_WIRE_1062;
wire	SYNTHESIZED_WIRE_1063;
wire	SYNTHESIZED_WIRE_1064;
wire	SYNTHESIZED_WIRE_1065;
wire	SYNTHESIZED_WIRE_1066;
wire	SYNTHESIZED_WIRE_1067;
wire	SYNTHESIZED_WIRE_1068;
wire	SYNTHESIZED_WIRE_1069;
wire	SYNTHESIZED_WIRE_1070;
wire	SYNTHESIZED_WIRE_1071;
wire	SYNTHESIZED_WIRE_1072;
wire	SYNTHESIZED_WIRE_1073;
wire	SYNTHESIZED_WIRE_1074;
wire	SYNTHESIZED_WIRE_1075;
wire	SYNTHESIZED_WIRE_1076;
wire	SYNTHESIZED_WIRE_1077;
wire	SYNTHESIZED_WIRE_1078;
wire	SYNTHESIZED_WIRE_1079;
wire	SYNTHESIZED_WIRE_1080;
wire	SYNTHESIZED_WIRE_1081;
wire	SYNTHESIZED_WIRE_1082;
wire	SYNTHESIZED_WIRE_1083;
wire	SYNTHESIZED_WIRE_1084;
wire	SYNTHESIZED_WIRE_1085;
wire	SYNTHESIZED_WIRE_1086;
wire	SYNTHESIZED_WIRE_1087;
wire	SYNTHESIZED_WIRE_1088;
wire	SYNTHESIZED_WIRE_1089;
wire	SYNTHESIZED_WIRE_1090;
wire	SYNTHESIZED_WIRE_1091;
wire	SYNTHESIZED_WIRE_1092;
wire	SYNTHESIZED_WIRE_1093;
wire	SYNTHESIZED_WIRE_1094;
wire	SYNTHESIZED_WIRE_1095;
wire	SYNTHESIZED_WIRE_1096;
wire	SYNTHESIZED_WIRE_1097;
wire	SYNTHESIZED_WIRE_1098;
wire	SYNTHESIZED_WIRE_1099;
wire	SYNTHESIZED_WIRE_1100;
wire	SYNTHESIZED_WIRE_1101;
wire	SYNTHESIZED_WIRE_1102;
wire	[47:0] SYNTHESIZED_WIRE_1103;





round	b2v_inst(
	.R1(SYNTHESIZED_WIRE_0),
	.R2(SYNTHESIZED_WIRE_1),
	.R3(SYNTHESIZED_WIRE_2),
	.R4(SYNTHESIZED_WIRE_3),
	.R5(SYNTHESIZED_WIRE_4),
	.R6(SYNTHESIZED_WIRE_5),
	.R7(SYNTHESIZED_WIRE_6),
	.R8(SYNTHESIZED_WIRE_7),
	.R9(SYNTHESIZED_WIRE_8),
	.R10(SYNTHESIZED_WIRE_9),
	.R11(SYNTHESIZED_WIRE_10),
	.R12(SYNTHESIZED_WIRE_11),
	.R13(SYNTHESIZED_WIRE_12),
	.R14(SYNTHESIZED_WIRE_13),
	.R15(SYNTHESIZED_WIRE_14),
	.R16(SYNTHESIZED_WIRE_15),
	.R17(SYNTHESIZED_WIRE_16),
	.R18(SYNTHESIZED_WIRE_17),
	.R19(SYNTHESIZED_WIRE_18),
	.R20(SYNTHESIZED_WIRE_19),
	.R21(SYNTHESIZED_WIRE_20),
	.R22(SYNTHESIZED_WIRE_21),
	.R23(SYNTHESIZED_WIRE_22),
	.R24(SYNTHESIZED_WIRE_23),
	.R25(SYNTHESIZED_WIRE_24),
	.R26(SYNTHESIZED_WIRE_25),
	.R27(SYNTHESIZED_WIRE_26),
	.R28(SYNTHESIZED_WIRE_27),
	.R29(SYNTHESIZED_WIRE_28),
	.R30(SYNTHESIZED_WIRE_29),
	.R31(SYNTHESIZED_WIRE_30),
	.R32(SYNTHESIZED_WIRE_31),
	.L1(SYNTHESIZED_WIRE_32),
	.L2(SYNTHESIZED_WIRE_33),
	.L3(SYNTHESIZED_WIRE_34),
	.L4(SYNTHESIZED_WIRE_35),
	.L5(SYNTHESIZED_WIRE_36),
	.L6(SYNTHESIZED_WIRE_37),
	.L7(SYNTHESIZED_WIRE_38),
	.L8(SYNTHESIZED_WIRE_39),
	.L9(SYNTHESIZED_WIRE_40),
	.L10(SYNTHESIZED_WIRE_41),
	.L11(SYNTHESIZED_WIRE_42),
	.L12(SYNTHESIZED_WIRE_43),
	.L13(SYNTHESIZED_WIRE_44),
	.L14(SYNTHESIZED_WIRE_45),
	.L15(SYNTHESIZED_WIRE_46),
	.L16(SYNTHESIZED_WIRE_47),
	.L17(SYNTHESIZED_WIRE_48),
	.L18(SYNTHESIZED_WIRE_49),
	.L19(SYNTHESIZED_WIRE_50),
	.L20(SYNTHESIZED_WIRE_51),
	.L21(SYNTHESIZED_WIRE_52),
	.L22(SYNTHESIZED_WIRE_53),
	.L23(SYNTHESIZED_WIRE_54),
	.L24(SYNTHESIZED_WIRE_55),
	.L25(SYNTHESIZED_WIRE_56),
	.L26(SYNTHESIZED_WIRE_57),
	.L27(SYNTHESIZED_WIRE_58),
	.L28(SYNTHESIZED_WIRE_59),
	.L29(SYNTHESIZED_WIRE_60),
	.L30(SYNTHESIZED_WIRE_61),
	.L31(SYNTHESIZED_WIRE_62),
	.L32(SYNTHESIZED_WIRE_63),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_64),
	.R_next1(SYNTHESIZED_WIRE_65),
	.R_next2(SYNTHESIZED_WIRE_66),
	.R_next3(SYNTHESIZED_WIRE_67),
	.R_next4(SYNTHESIZED_WIRE_68),
	.R_next5(SYNTHESIZED_WIRE_69),
	.R_next6(SYNTHESIZED_WIRE_70),
	.R_next7(SYNTHESIZED_WIRE_71),
	.R_next8(SYNTHESIZED_WIRE_72),
	.R_next9(SYNTHESIZED_WIRE_73),
	.R_next10(SYNTHESIZED_WIRE_74),
	.R_next11(SYNTHESIZED_WIRE_75),
	.R_next12(SYNTHESIZED_WIRE_76),
	.R_next13(SYNTHESIZED_WIRE_77),
	.R_next14(SYNTHESIZED_WIRE_78),
	.R_next15(SYNTHESIZED_WIRE_79),
	.R_next16(SYNTHESIZED_WIRE_80),
	.R_next17(SYNTHESIZED_WIRE_81),
	.R_next18(SYNTHESIZED_WIRE_82),
	.R_next19(SYNTHESIZED_WIRE_83),
	.R_next20(SYNTHESIZED_WIRE_84),
	.R_next21(SYNTHESIZED_WIRE_85),
	.R_next22(SYNTHESIZED_WIRE_86),
	.R_next23(SYNTHESIZED_WIRE_87),
	.R_next24(SYNTHESIZED_WIRE_88),
	.R_next25(SYNTHESIZED_WIRE_89),
	.R_next26(SYNTHESIZED_WIRE_90),
	.R_next27(SYNTHESIZED_WIRE_91),
	.R_next28(SYNTHESIZED_WIRE_92),
	.R_next29(SYNTHESIZED_WIRE_93),
	.R_next30(SYNTHESIZED_WIRE_94),
	.R_next31(SYNTHESIZED_WIRE_95),
	.R_next32(SYNTHESIZED_WIRE_96),
	.L_next1(SYNTHESIZED_WIRE_97),
	.L_next2(SYNTHESIZED_WIRE_98),
	.L_next3(SYNTHESIZED_WIRE_99),
	.L_next4(SYNTHESIZED_WIRE_100),
	.L_next5(SYNTHESIZED_WIRE_101),
	.L_next6(SYNTHESIZED_WIRE_102),
	.L_next7(SYNTHESIZED_WIRE_103),
	.L_next8(SYNTHESIZED_WIRE_104),
	.L_next9(SYNTHESIZED_WIRE_105),
	.L_next10(SYNTHESIZED_WIRE_106),
	.L_next11(SYNTHESIZED_WIRE_107),
	.L_next12(SYNTHESIZED_WIRE_108),
	.L_next13(SYNTHESIZED_WIRE_109),
	.L_next14(SYNTHESIZED_WIRE_110),
	.L_next15(SYNTHESIZED_WIRE_111),
	.L_next16(SYNTHESIZED_WIRE_112),
	.L_next17(SYNTHESIZED_WIRE_113),
	.L_next18(SYNTHESIZED_WIRE_114),
	.L_next19(SYNTHESIZED_WIRE_115),
	.L_next20(SYNTHESIZED_WIRE_116),
	.L_next21(SYNTHESIZED_WIRE_117),
	.L_next22(SYNTHESIZED_WIRE_118),
	.L_next23(SYNTHESIZED_WIRE_119),
	.L_next24(SYNTHESIZED_WIRE_120),
	.L_next25(SYNTHESIZED_WIRE_121),
	.L_next26(SYNTHESIZED_WIRE_122),
	.L_next27(SYNTHESIZED_WIRE_123),
	.L_next28(SYNTHESIZED_WIRE_124),
	.L_next29(SYNTHESIZED_WIRE_125),
	.L_next30(SYNTHESIZED_WIRE_126),
	.L_next31(SYNTHESIZED_WIRE_127),
	.L_next32(SYNTHESIZED_WIRE_128));


key_generator	b2v_inst1(
	.initial_key(initial_key),
	.round10key(SYNTHESIZED_WIRE_713),
	.round11key(SYNTHESIZED_WIRE_778),
	.round12key(SYNTHESIZED_WIRE_843),
	.round13key(SYNTHESIZED_WIRE_908),
	.round14key(SYNTHESIZED_WIRE_973),
	.round15key(SYNTHESIZED_WIRE_1038),
	.round16key(SYNTHESIZED_WIRE_1103),
	.round1key(SYNTHESIZED_WIRE_64),
	.round2key(SYNTHESIZED_WIRE_129),
	.round3key(SYNTHESIZED_WIRE_194),
	.round4key(SYNTHESIZED_WIRE_323),
	.round5key(SYNTHESIZED_WIRE_388),
	.round6key(SYNTHESIZED_WIRE_453),
	.round7key(SYNTHESIZED_WIRE_518),
	.round8key(SYNTHESIZED_WIRE_583),
	.round9key(SYNTHESIZED_WIRE_648));


IP	b2v_inst3(
	.ip_in1(reg10),
	.ip_in2(reg11),
	.ip_in3(reg12),
	.ip_in4(reg13),
	.ip_in5(reg2[0]),
	.ip_in6(reg2[1]),
	.ip_in7(reg2[2]),
	.ip_in8(reg2[3]),
	.ip_in9(reg3[0]),
	.ip_in10(reg3[1]),
	.ip_in11(reg3[2]),
	.ip_in12(reg3[3]),
	.ip_in13(reg4[0]),
	.ip_in14(reg4[1]),
	.ip_in15(reg4[2]),
	.ip_in16(reg4[3]),
	.ip_in17(reg5[0]),
	.ip_in18(reg5[1]),
	.ip_in19(reg5[2]),
	.ip_in20(reg5[3]),
	.ip_in21(reg6[0]),
	.ip_in22(reg6[1]),
	.ip_in23(reg6[2]),
	.ip_in24(reg6[3]),
	.ip_in25(reg7[0]),
	.ip_in26(reg7[1]),
	.ip_in27(reg7[2]),
	.ip_in28(reg7[3]),
	.ip_in29(reg8[0]),
	.ip_in30(reg8[1]),
	.ip_in31(reg8[2]),
	.ip_in32(reg8[3]),
	.ip_in33(reg9[0]),
	.ip_in34(reg9[1]),
	.ip_in35(reg9[2]),
	.ip_in36(reg9[3]),
	.ip_in37(reg100),
	.ip_in38(reg101),
	.ip_in39(reg102),
	.ip_in40(reg103),
	.ip_in41(reg110),
	.ip_in42(reg111),
	.ip_in43(reg112),
	.ip_in44(reg113),
	.ip_in45(reg120),
	.ip_in46(reg121),
	.ip_in47(reg122),
	.ip_in48(reg123),
	.ip_in49(reg130),
	.ip_in50(reg131),
	.ip_in51(reg132),
	.ip_in52(reg133),
	.ip_in53(reg14[0]),
	.ip_in54(reg14[1]),
	.ip_in55(reg14[2]),
	.ip_in56(reg14[3]),
	.ip_in57(reg15[0]),
	.ip_in58(reg15[1]),
	.ip_in59(reg15[2]),
	.ip_in60(reg15[3]),
	.ip_in61(reg16[0]),
	.ip_in62(reg16[1]),
	.ip_in63(reg16[2]),
	.ip_in64(reg16[3]),
	.ip_out1(SYNTHESIZED_WIRE_0),
	.ip_out2(SYNTHESIZED_WIRE_1),
	.ip_out3(SYNTHESIZED_WIRE_2),
	.ip_out4(SYNTHESIZED_WIRE_3),
	.ip_out5(SYNTHESIZED_WIRE_4),
	.ip_out6(SYNTHESIZED_WIRE_5),
	.ip_out7(SYNTHESIZED_WIRE_6),
	.ip_out8(SYNTHESIZED_WIRE_7),
	.ip_out9(SYNTHESIZED_WIRE_8),
	.ip_out10(SYNTHESIZED_WIRE_9),
	.ip_out11(SYNTHESIZED_WIRE_10),
	.ip_out12(SYNTHESIZED_WIRE_11),
	.ip_out13(SYNTHESIZED_WIRE_12),
	.ip_out14(SYNTHESIZED_WIRE_13),
	.ip_out15(SYNTHESIZED_WIRE_14),
	.ip_out16(SYNTHESIZED_WIRE_15),
	.ip_out17(SYNTHESIZED_WIRE_16),
	.ip_out18(SYNTHESIZED_WIRE_17),
	.ip_out19(SYNTHESIZED_WIRE_18),
	.ip_out20(SYNTHESIZED_WIRE_19),
	.ip_out21(SYNTHESIZED_WIRE_20),
	.ip_out22(SYNTHESIZED_WIRE_21),
	.ip_out23(SYNTHESIZED_WIRE_22),
	.ip_out24(SYNTHESIZED_WIRE_23),
	.ip_out25(SYNTHESIZED_WIRE_24),
	.ip_out26(SYNTHESIZED_WIRE_25),
	.ip_out27(SYNTHESIZED_WIRE_26),
	.ip_out28(SYNTHESIZED_WIRE_27),
	.ip_out29(SYNTHESIZED_WIRE_28),
	.ip_out30(SYNTHESIZED_WIRE_29),
	.ip_out31(SYNTHESIZED_WIRE_30),
	.ip_out32(SYNTHESIZED_WIRE_31),
	.ip_out33(SYNTHESIZED_WIRE_32),
	.ip_out34(SYNTHESIZED_WIRE_33),
	.ip_out35(SYNTHESIZED_WIRE_34),
	.ip_out36(SYNTHESIZED_WIRE_35),
	.ip_out37(SYNTHESIZED_WIRE_36),
	.ip_out38(SYNTHESIZED_WIRE_37),
	.ip_out39(SYNTHESIZED_WIRE_38),
	.ip_out40(SYNTHESIZED_WIRE_39),
	.ip_out41(SYNTHESIZED_WIRE_40),
	.ip_out42(SYNTHESIZED_WIRE_41),
	.ip_out43(SYNTHESIZED_WIRE_42),
	.ip_out44(SYNTHESIZED_WIRE_43),
	.ip_out45(SYNTHESIZED_WIRE_44),
	.ip_out46(SYNTHESIZED_WIRE_45),
	.ip_out47(SYNTHESIZED_WIRE_46),
	.ip_out48(SYNTHESIZED_WIRE_47),
	.ip_out49(SYNTHESIZED_WIRE_48),
	.ip_out50(SYNTHESIZED_WIRE_49),
	.ip_out51(SYNTHESIZED_WIRE_50),
	.ip_out52(SYNTHESIZED_WIRE_51),
	.ip_out53(SYNTHESIZED_WIRE_52),
	.ip_out54(SYNTHESIZED_WIRE_53),
	.ip_out55(SYNTHESIZED_WIRE_54),
	.ip_out56(SYNTHESIZED_WIRE_55),
	.ip_out57(SYNTHESIZED_WIRE_56),
	.ip_out58(SYNTHESIZED_WIRE_57),
	.ip_out59(SYNTHESIZED_WIRE_58),
	.ip_out60(SYNTHESIZED_WIRE_59),
	.ip_out61(SYNTHESIZED_WIRE_60),
	.ip_out62(SYNTHESIZED_WIRE_61),
	.ip_out63(SYNTHESIZED_WIRE_62),
	.ip_out64(SYNTHESIZED_WIRE_63));


round	b2v_inst41(
	.R1(SYNTHESIZED_WIRE_65),
	.R2(SYNTHESIZED_WIRE_66),
	.R3(SYNTHESIZED_WIRE_67),
	.R4(SYNTHESIZED_WIRE_68),
	.R5(SYNTHESIZED_WIRE_69),
	.R6(SYNTHESIZED_WIRE_70),
	.R7(SYNTHESIZED_WIRE_71),
	.R8(SYNTHESIZED_WIRE_72),
	.R9(SYNTHESIZED_WIRE_73),
	.R10(SYNTHESIZED_WIRE_74),
	.R11(SYNTHESIZED_WIRE_75),
	.R12(SYNTHESIZED_WIRE_76),
	.R13(SYNTHESIZED_WIRE_77),
	.R14(SYNTHESIZED_WIRE_78),
	.R15(SYNTHESIZED_WIRE_79),
	.R16(SYNTHESIZED_WIRE_80),
	.R17(SYNTHESIZED_WIRE_81),
	.R18(SYNTHESIZED_WIRE_82),
	.R19(SYNTHESIZED_WIRE_83),
	.R20(SYNTHESIZED_WIRE_84),
	.R21(SYNTHESIZED_WIRE_85),
	.R22(SYNTHESIZED_WIRE_86),
	.R23(SYNTHESIZED_WIRE_87),
	.R24(SYNTHESIZED_WIRE_88),
	.R25(SYNTHESIZED_WIRE_89),
	.R26(SYNTHESIZED_WIRE_90),
	.R27(SYNTHESIZED_WIRE_91),
	.R28(SYNTHESIZED_WIRE_92),
	.R29(SYNTHESIZED_WIRE_93),
	.R30(SYNTHESIZED_WIRE_94),
	.R31(SYNTHESIZED_WIRE_95),
	.R32(SYNTHESIZED_WIRE_96),
	.L1(SYNTHESIZED_WIRE_97),
	.L2(SYNTHESIZED_WIRE_98),
	.L3(SYNTHESIZED_WIRE_99),
	.L4(SYNTHESIZED_WIRE_100),
	.L5(SYNTHESIZED_WIRE_101),
	.L6(SYNTHESIZED_WIRE_102),
	.L7(SYNTHESIZED_WIRE_103),
	.L8(SYNTHESIZED_WIRE_104),
	.L9(SYNTHESIZED_WIRE_105),
	.L10(SYNTHESIZED_WIRE_106),
	.L11(SYNTHESIZED_WIRE_107),
	.L12(SYNTHESIZED_WIRE_108),
	.L13(SYNTHESIZED_WIRE_109),
	.L14(SYNTHESIZED_WIRE_110),
	.L15(SYNTHESIZED_WIRE_111),
	.L16(SYNTHESIZED_WIRE_112),
	.L17(SYNTHESIZED_WIRE_113),
	.L18(SYNTHESIZED_WIRE_114),
	.L19(SYNTHESIZED_WIRE_115),
	.L20(SYNTHESIZED_WIRE_116),
	.L21(SYNTHESIZED_WIRE_117),
	.L22(SYNTHESIZED_WIRE_118),
	.L23(SYNTHESIZED_WIRE_119),
	.L24(SYNTHESIZED_WIRE_120),
	.L25(SYNTHESIZED_WIRE_121),
	.L26(SYNTHESIZED_WIRE_122),
	.L27(SYNTHESIZED_WIRE_123),
	.L28(SYNTHESIZED_WIRE_124),
	.L29(SYNTHESIZED_WIRE_125),
	.L30(SYNTHESIZED_WIRE_126),
	.L31(SYNTHESIZED_WIRE_127),
	.L32(SYNTHESIZED_WIRE_128),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_129),
	.R_next1(SYNTHESIZED_WIRE_130),
	.R_next2(SYNTHESIZED_WIRE_131),
	.R_next3(SYNTHESIZED_WIRE_132),
	.R_next4(SYNTHESIZED_WIRE_133),
	.R_next5(SYNTHESIZED_WIRE_134),
	.R_next6(SYNTHESIZED_WIRE_135),
	.R_next7(SYNTHESIZED_WIRE_136),
	.R_next8(SYNTHESIZED_WIRE_137),
	.R_next9(SYNTHESIZED_WIRE_138),
	.R_next10(SYNTHESIZED_WIRE_139),
	.R_next11(SYNTHESIZED_WIRE_140),
	.R_next12(SYNTHESIZED_WIRE_141),
	.R_next13(SYNTHESIZED_WIRE_142),
	.R_next14(SYNTHESIZED_WIRE_143),
	.R_next15(SYNTHESIZED_WIRE_144),
	.R_next16(SYNTHESIZED_WIRE_145),
	.R_next17(SYNTHESIZED_WIRE_146),
	.R_next18(SYNTHESIZED_WIRE_147),
	.R_next19(SYNTHESIZED_WIRE_148),
	.R_next20(SYNTHESIZED_WIRE_149),
	.R_next21(SYNTHESIZED_WIRE_150),
	.R_next22(SYNTHESIZED_WIRE_151),
	.R_next23(SYNTHESIZED_WIRE_152),
	.R_next24(SYNTHESIZED_WIRE_153),
	.R_next25(SYNTHESIZED_WIRE_154),
	.R_next26(SYNTHESIZED_WIRE_155),
	.R_next27(SYNTHESIZED_WIRE_156),
	.R_next28(SYNTHESIZED_WIRE_157),
	.R_next29(SYNTHESIZED_WIRE_158),
	.R_next30(SYNTHESIZED_WIRE_159),
	.R_next31(SYNTHESIZED_WIRE_160),
	.R_next32(SYNTHESIZED_WIRE_161),
	.L_next1(SYNTHESIZED_WIRE_162),
	.L_next2(SYNTHESIZED_WIRE_163),
	.L_next3(SYNTHESIZED_WIRE_164),
	.L_next4(SYNTHESIZED_WIRE_165),
	.L_next5(SYNTHESIZED_WIRE_166),
	.L_next6(SYNTHESIZED_WIRE_167),
	.L_next7(SYNTHESIZED_WIRE_168),
	.L_next8(SYNTHESIZED_WIRE_169),
	.L_next9(SYNTHESIZED_WIRE_170),
	.L_next10(SYNTHESIZED_WIRE_171),
	.L_next11(SYNTHESIZED_WIRE_172),
	.L_next12(SYNTHESIZED_WIRE_173),
	.L_next13(SYNTHESIZED_WIRE_174),
	.L_next14(SYNTHESIZED_WIRE_175),
	.L_next15(SYNTHESIZED_WIRE_176),
	.L_next16(SYNTHESIZED_WIRE_177),
	.L_next17(SYNTHESIZED_WIRE_178),
	.L_next18(SYNTHESIZED_WIRE_179),
	.L_next19(SYNTHESIZED_WIRE_180),
	.L_next20(SYNTHESIZED_WIRE_181),
	.L_next21(SYNTHESIZED_WIRE_182),
	.L_next22(SYNTHESIZED_WIRE_183),
	.L_next23(SYNTHESIZED_WIRE_184),
	.L_next24(SYNTHESIZED_WIRE_185),
	.L_next25(SYNTHESIZED_WIRE_186),
	.L_next26(SYNTHESIZED_WIRE_187),
	.L_next27(SYNTHESIZED_WIRE_188),
	.L_next28(SYNTHESIZED_WIRE_189),
	.L_next29(SYNTHESIZED_WIRE_190),
	.L_next30(SYNTHESIZED_WIRE_191),
	.L_next31(SYNTHESIZED_WIRE_192),
	.L_next32(SYNTHESIZED_WIRE_193));


round	b2v_inst42(
	.R1(SYNTHESIZED_WIRE_130),
	.R2(SYNTHESIZED_WIRE_131),
	.R3(SYNTHESIZED_WIRE_132),
	.R4(SYNTHESIZED_WIRE_133),
	.R5(SYNTHESIZED_WIRE_134),
	.R6(SYNTHESIZED_WIRE_135),
	.R7(SYNTHESIZED_WIRE_136),
	.R8(SYNTHESIZED_WIRE_137),
	.R9(SYNTHESIZED_WIRE_138),
	.R10(SYNTHESIZED_WIRE_139),
	.R11(SYNTHESIZED_WIRE_140),
	.R12(SYNTHESIZED_WIRE_141),
	.R13(SYNTHESIZED_WIRE_142),
	.R14(SYNTHESIZED_WIRE_143),
	.R15(SYNTHESIZED_WIRE_144),
	.R16(SYNTHESIZED_WIRE_145),
	.R17(SYNTHESIZED_WIRE_146),
	.R18(SYNTHESIZED_WIRE_147),
	.R19(SYNTHESIZED_WIRE_148),
	.R20(SYNTHESIZED_WIRE_149),
	.R21(SYNTHESIZED_WIRE_150),
	.R22(SYNTHESIZED_WIRE_151),
	.R23(SYNTHESIZED_WIRE_152),
	.R24(SYNTHESIZED_WIRE_153),
	.R25(SYNTHESIZED_WIRE_154),
	.R26(SYNTHESIZED_WIRE_155),
	.R27(SYNTHESIZED_WIRE_156),
	.R28(SYNTHESIZED_WIRE_157),
	.R29(SYNTHESIZED_WIRE_158),
	.R30(SYNTHESIZED_WIRE_159),
	.R31(SYNTHESIZED_WIRE_160),
	.R32(SYNTHESIZED_WIRE_161),
	.L1(SYNTHESIZED_WIRE_162),
	.L2(SYNTHESIZED_WIRE_163),
	.L3(SYNTHESIZED_WIRE_164),
	.L4(SYNTHESIZED_WIRE_165),
	.L5(SYNTHESIZED_WIRE_166),
	.L6(SYNTHESIZED_WIRE_167),
	.L7(SYNTHESIZED_WIRE_168),
	.L8(SYNTHESIZED_WIRE_169),
	.L9(SYNTHESIZED_WIRE_170),
	.L10(SYNTHESIZED_WIRE_171),
	.L11(SYNTHESIZED_WIRE_172),
	.L12(SYNTHESIZED_WIRE_173),
	.L13(SYNTHESIZED_WIRE_174),
	.L14(SYNTHESIZED_WIRE_175),
	.L15(SYNTHESIZED_WIRE_176),
	.L16(SYNTHESIZED_WIRE_177),
	.L17(SYNTHESIZED_WIRE_178),
	.L18(SYNTHESIZED_WIRE_179),
	.L19(SYNTHESIZED_WIRE_180),
	.L20(SYNTHESIZED_WIRE_181),
	.L21(SYNTHESIZED_WIRE_182),
	.L22(SYNTHESIZED_WIRE_183),
	.L23(SYNTHESIZED_WIRE_184),
	.L24(SYNTHESIZED_WIRE_185),
	.L25(SYNTHESIZED_WIRE_186),
	.L26(SYNTHESIZED_WIRE_187),
	.L27(SYNTHESIZED_WIRE_188),
	.L28(SYNTHESIZED_WIRE_189),
	.L29(SYNTHESIZED_WIRE_190),
	.L30(SYNTHESIZED_WIRE_191),
	.L31(SYNTHESIZED_WIRE_192),
	.L32(SYNTHESIZED_WIRE_193),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_194),
	.R_next1(SYNTHESIZED_WIRE_259),
	.R_next2(SYNTHESIZED_WIRE_260),
	.R_next3(SYNTHESIZED_WIRE_261),
	.R_next4(SYNTHESIZED_WIRE_262),
	.R_next5(SYNTHESIZED_WIRE_263),
	.R_next6(SYNTHESIZED_WIRE_264),
	.R_next7(SYNTHESIZED_WIRE_265),
	.R_next8(SYNTHESIZED_WIRE_266),
	.R_next9(SYNTHESIZED_WIRE_267),
	.R_next10(SYNTHESIZED_WIRE_268),
	.R_next11(SYNTHESIZED_WIRE_269),
	.R_next12(SYNTHESIZED_WIRE_270),
	.R_next13(SYNTHESIZED_WIRE_271),
	.R_next14(SYNTHESIZED_WIRE_272),
	.R_next15(SYNTHESIZED_WIRE_273),
	.R_next16(SYNTHESIZED_WIRE_274),
	.R_next17(SYNTHESIZED_WIRE_275),
	.R_next18(SYNTHESIZED_WIRE_276),
	.R_next19(SYNTHESIZED_WIRE_277),
	.R_next20(SYNTHESIZED_WIRE_278),
	.R_next21(SYNTHESIZED_WIRE_279),
	.R_next22(SYNTHESIZED_WIRE_280),
	.R_next23(SYNTHESIZED_WIRE_281),
	.R_next24(SYNTHESIZED_WIRE_282),
	.R_next25(SYNTHESIZED_WIRE_283),
	.R_next26(SYNTHESIZED_WIRE_284),
	.R_next27(SYNTHESIZED_WIRE_285),
	.R_next28(SYNTHESIZED_WIRE_286),
	.R_next29(SYNTHESIZED_WIRE_287),
	.R_next30(SYNTHESIZED_WIRE_288),
	.R_next31(SYNTHESIZED_WIRE_289),
	.R_next32(SYNTHESIZED_WIRE_290),
	.L_next1(SYNTHESIZED_WIRE_291),
	.L_next2(SYNTHESIZED_WIRE_292),
	.L_next3(SYNTHESIZED_WIRE_293),
	.L_next4(SYNTHESIZED_WIRE_294),
	.L_next5(SYNTHESIZED_WIRE_295),
	.L_next6(SYNTHESIZED_WIRE_296),
	.L_next7(SYNTHESIZED_WIRE_297),
	.L_next8(SYNTHESIZED_WIRE_298),
	.L_next9(SYNTHESIZED_WIRE_299),
	.L_next10(SYNTHESIZED_WIRE_300),
	.L_next11(SYNTHESIZED_WIRE_301),
	.L_next12(SYNTHESIZED_WIRE_302),
	.L_next13(SYNTHESIZED_WIRE_303),
	.L_next14(SYNTHESIZED_WIRE_304),
	.L_next15(SYNTHESIZED_WIRE_305),
	.L_next16(SYNTHESIZED_WIRE_306),
	.L_next17(SYNTHESIZED_WIRE_307),
	.L_next18(SYNTHESIZED_WIRE_308),
	.L_next19(SYNTHESIZED_WIRE_309),
	.L_next20(SYNTHESIZED_WIRE_310),
	.L_next21(SYNTHESIZED_WIRE_311),
	.L_next22(SYNTHESIZED_WIRE_312),
	.L_next23(SYNTHESIZED_WIRE_313),
	.L_next24(SYNTHESIZED_WIRE_314),
	.L_next25(SYNTHESIZED_WIRE_315),
	.L_next26(SYNTHESIZED_WIRE_316),
	.L_next27(SYNTHESIZED_WIRE_317),
	.L_next28(SYNTHESIZED_WIRE_318),
	.L_next29(SYNTHESIZED_WIRE_319),
	.L_next30(SYNTHESIZED_WIRE_320),
	.L_next31(SYNTHESIZED_WIRE_321),
	.L_next32(SYNTHESIZED_WIRE_322));


IP_inv	b2v_inst43(
	.ipinv_in1(SYNTHESIZED_WIRE_195),
	.ipinv_in2(SYNTHESIZED_WIRE_196),
	.ipinv_in3(SYNTHESIZED_WIRE_197),
	.ipinv_in4(SYNTHESIZED_WIRE_198),
	.ipinv_in5(SYNTHESIZED_WIRE_199),
	.ipinv_in6(SYNTHESIZED_WIRE_200),
	.ipinv_in7(SYNTHESIZED_WIRE_201),
	.ipinv_in8(SYNTHESIZED_WIRE_202),
	.ipinv_in9(SYNTHESIZED_WIRE_203),
	.ipinv_in10(SYNTHESIZED_WIRE_204),
	.ipinv_in11(SYNTHESIZED_WIRE_205),
	.ipinv_in12(SYNTHESIZED_WIRE_206),
	.ipinv_in13(SYNTHESIZED_WIRE_207),
	.ipinv_in14(SYNTHESIZED_WIRE_208),
	.ipinv_in15(SYNTHESIZED_WIRE_209),
	.ipinv_in16(SYNTHESIZED_WIRE_210),
	.ipinv_in17(SYNTHESIZED_WIRE_211),
	.ipinv_in18(SYNTHESIZED_WIRE_212),
	.ipinv_in19(SYNTHESIZED_WIRE_213),
	.ipinv_in20(SYNTHESIZED_WIRE_214),
	.ipinv_in21(SYNTHESIZED_WIRE_215),
	.ipinv_in22(SYNTHESIZED_WIRE_216),
	.ipinv_in23(SYNTHESIZED_WIRE_217),
	.ipinv_in24(SYNTHESIZED_WIRE_218),
	.ipinv_in25(SYNTHESIZED_WIRE_219),
	.ipinv_in26(SYNTHESIZED_WIRE_220),
	.ipinv_in27(SYNTHESIZED_WIRE_221),
	.ipinv_in28(SYNTHESIZED_WIRE_222),
	.ipinv_in29(SYNTHESIZED_WIRE_223),
	.ipinv_in30(SYNTHESIZED_WIRE_224),
	.ipinv_in31(SYNTHESIZED_WIRE_225),
	.ipinv_in32(SYNTHESIZED_WIRE_226),
	.ipinv_in33(SYNTHESIZED_WIRE_227),
	.ipinv_in34(SYNTHESIZED_WIRE_228),
	.ipinv_in35(SYNTHESIZED_WIRE_229),
	.ipinv_in36(SYNTHESIZED_WIRE_230),
	.ipinv_in37(SYNTHESIZED_WIRE_231),
	.ipinv_in38(SYNTHESIZED_WIRE_232),
	.ipinv_in39(SYNTHESIZED_WIRE_233),
	.ipinv_in40(SYNTHESIZED_WIRE_234),
	.ipinv_in41(SYNTHESIZED_WIRE_235),
	.ipinv_in42(SYNTHESIZED_WIRE_236),
	.ipinv_in43(SYNTHESIZED_WIRE_237),
	.ipinv_in44(SYNTHESIZED_WIRE_238),
	.ipinv_in45(SYNTHESIZED_WIRE_239),
	.ipinv_in46(SYNTHESIZED_WIRE_240),
	.ipinv_in47(SYNTHESIZED_WIRE_241),
	.ipinv_in48(SYNTHESIZED_WIRE_242),
	.ipinv_in49(SYNTHESIZED_WIRE_243),
	.ipinv_in50(SYNTHESIZED_WIRE_244),
	.ipinv_in51(SYNTHESIZED_WIRE_245),
	.ipinv_in52(SYNTHESIZED_WIRE_246),
	.ipinv_in53(SYNTHESIZED_WIRE_247),
	.ipinv_in54(SYNTHESIZED_WIRE_248),
	.ipinv_in55(SYNTHESIZED_WIRE_249),
	.ipinv_in56(SYNTHESIZED_WIRE_250),
	.ipinv_in57(SYNTHESIZED_WIRE_251),
	.ipinv_in58(SYNTHESIZED_WIRE_252),
	.ipinv_in59(SYNTHESIZED_WIRE_253),
	.ipinv_in60(SYNTHESIZED_WIRE_254),
	.ipinv_in61(SYNTHESIZED_WIRE_255),
	.ipinv_in62(SYNTHESIZED_WIRE_256),
	.ipinv_in63(SYNTHESIZED_WIRE_257),
	.ipinv_in64(SYNTHESIZED_WIRE_258),
	.ipinv_out1(des_encrypt_out_ALTERA_SYNTHESIZED[0]),
	.ipinv_out2(des_encrypt_out_ALTERA_SYNTHESIZED[1]),
	.ipinv_out3(des_encrypt_out_ALTERA_SYNTHESIZED[2]),
	.ipinv_out4(des_encrypt_out_ALTERA_SYNTHESIZED[3]),
	.ipinv_out5(des_encrypt_out_ALTERA_SYNTHESIZED[4]),
	.ipinv_out6(des_encrypt_out_ALTERA_SYNTHESIZED[5]),
	.ipinv_out7(des_encrypt_out_ALTERA_SYNTHESIZED[6]),
	.ipinv_out8(des_encrypt_out_ALTERA_SYNTHESIZED[7]),
	.ipinv_out9(des_encrypt_out_ALTERA_SYNTHESIZED[8]),
	.ipinv_out10(des_encrypt_out_ALTERA_SYNTHESIZED[9]),
	.ipinv_out11(des_encrypt_out_ALTERA_SYNTHESIZED[10]),
	.ipinv_out12(des_encrypt_out_ALTERA_SYNTHESIZED[11]),
	.ipinv_out13(des_encrypt_out_ALTERA_SYNTHESIZED[12]),
	.ipinv_out14(des_encrypt_out_ALTERA_SYNTHESIZED[13]),
	.ipinv_out15(des_encrypt_out_ALTERA_SYNTHESIZED[14]),
	.ipinv_out16(des_encrypt_out_ALTERA_SYNTHESIZED[15]),
	.ipinv_out17(des_encrypt_out_ALTERA_SYNTHESIZED[16]),
	.ipinv_out18(des_encrypt_out_ALTERA_SYNTHESIZED[17]),
	.ipinv_out19(des_encrypt_out_ALTERA_SYNTHESIZED[18]),
	.ipinv_out20(des_encrypt_out_ALTERA_SYNTHESIZED[19]),
	.ipinv_out21(des_encrypt_out_ALTERA_SYNTHESIZED[20]),
	.ipinv_out22(des_encrypt_out_ALTERA_SYNTHESIZED[21]),
	.ipinv_out23(des_encrypt_out_ALTERA_SYNTHESIZED[22]),
	.ipinv_out24(des_encrypt_out_ALTERA_SYNTHESIZED[23]),
	.ipinv_out25(des_encrypt_out_ALTERA_SYNTHESIZED[24]),
	.ipinv_out26(des_encrypt_out_ALTERA_SYNTHESIZED[25]),
	.ipinv_out27(des_encrypt_out_ALTERA_SYNTHESIZED[26]),
	.ipinv_out28(des_encrypt_out_ALTERA_SYNTHESIZED[27]),
	.ipinv_out29(des_encrypt_out_ALTERA_SYNTHESIZED[28]),
	.ipinv_out30(des_encrypt_out_ALTERA_SYNTHESIZED[29]),
	.ipinv_out31(des_encrypt_out_ALTERA_SYNTHESIZED[30]),
	.ipinv_out32(des_encrypt_out_ALTERA_SYNTHESIZED[31]),
	.ipinv_out33(des_encrypt_out_ALTERA_SYNTHESIZED[32]),
	.ipinv_out34(des_encrypt_out_ALTERA_SYNTHESIZED[33]),
	.ipinv_out35(des_encrypt_out_ALTERA_SYNTHESIZED[34]),
	.ipinv_out36(des_encrypt_out_ALTERA_SYNTHESIZED[35]),
	.ipinv_out37(des_encrypt_out_ALTERA_SYNTHESIZED[36]),
	.ipinv_out38(des_encrypt_out_ALTERA_SYNTHESIZED[37]),
	.ipinv_out39(des_encrypt_out_ALTERA_SYNTHESIZED[38]),
	.ipinv_out40(des_encrypt_out_ALTERA_SYNTHESIZED[39]),
	.ipinv_out41(des_encrypt_out_ALTERA_SYNTHESIZED[40]),
	.ipinv_out42(des_encrypt_out_ALTERA_SYNTHESIZED[41]),
	.ipinv_out43(des_encrypt_out_ALTERA_SYNTHESIZED[42]),
	.ipinv_out44(des_encrypt_out_ALTERA_SYNTHESIZED[43]),
	.ipinv_out45(des_encrypt_out_ALTERA_SYNTHESIZED[44]),
	.ipinv_out46(des_encrypt_out_ALTERA_SYNTHESIZED[45]),
	.ipinv_out47(des_encrypt_out_ALTERA_SYNTHESIZED[46]),
	.ipinv_out48(des_encrypt_out_ALTERA_SYNTHESIZED[47]),
	.ipinv_out49(des_encrypt_out_ALTERA_SYNTHESIZED[48]),
	.ipinv_out50(des_encrypt_out_ALTERA_SYNTHESIZED[49]),
	.ipinv_out51(des_encrypt_out_ALTERA_SYNTHESIZED[50]),
	.ipinv_out52(des_encrypt_out_ALTERA_SYNTHESIZED[51]),
	.ipinv_out53(des_encrypt_out_ALTERA_SYNTHESIZED[52]),
	.ipinv_out54(des_encrypt_out_ALTERA_SYNTHESIZED[53]),
	.ipinv_out55(des_encrypt_out_ALTERA_SYNTHESIZED[54]),
	.ipinv_out56(des_encrypt_out_ALTERA_SYNTHESIZED[55]),
	.ipinv_out57(des_encrypt_out_ALTERA_SYNTHESIZED[56]),
	.ipinv_out58(des_encrypt_out_ALTERA_SYNTHESIZED[57]),
	.ipinv_out59(des_encrypt_out_ALTERA_SYNTHESIZED[58]),
	.ipinv_out60(des_encrypt_out_ALTERA_SYNTHESIZED[59]),
	.ipinv_out61(des_encrypt_out_ALTERA_SYNTHESIZED[60]),
	.ipinv_out62(des_encrypt_out_ALTERA_SYNTHESIZED[61]),
	.ipinv_out63(des_encrypt_out_ALTERA_SYNTHESIZED[62]),
	.ipinv_out64(des_encrypt_out_ALTERA_SYNTHESIZED[63]));


round	b2v_inst431(
	.R1(SYNTHESIZED_WIRE_259),
	.R2(SYNTHESIZED_WIRE_260),
	.R3(SYNTHESIZED_WIRE_261),
	.R4(SYNTHESIZED_WIRE_262),
	.R5(SYNTHESIZED_WIRE_263),
	.R6(SYNTHESIZED_WIRE_264),
	.R7(SYNTHESIZED_WIRE_265),
	.R8(SYNTHESIZED_WIRE_266),
	.R9(SYNTHESIZED_WIRE_267),
	.R10(SYNTHESIZED_WIRE_268),
	.R11(SYNTHESIZED_WIRE_269),
	.R12(SYNTHESIZED_WIRE_270),
	.R13(SYNTHESIZED_WIRE_271),
	.R14(SYNTHESIZED_WIRE_272),
	.R15(SYNTHESIZED_WIRE_273),
	.R16(SYNTHESIZED_WIRE_274),
	.R17(SYNTHESIZED_WIRE_275),
	.R18(SYNTHESIZED_WIRE_276),
	.R19(SYNTHESIZED_WIRE_277),
	.R20(SYNTHESIZED_WIRE_278),
	.R21(SYNTHESIZED_WIRE_279),
	.R22(SYNTHESIZED_WIRE_280),
	.R23(SYNTHESIZED_WIRE_281),
	.R24(SYNTHESIZED_WIRE_282),
	.R25(SYNTHESIZED_WIRE_283),
	.R26(SYNTHESIZED_WIRE_284),
	.R27(SYNTHESIZED_WIRE_285),
	.R28(SYNTHESIZED_WIRE_286),
	.R29(SYNTHESIZED_WIRE_287),
	.R30(SYNTHESIZED_WIRE_288),
	.R31(SYNTHESIZED_WIRE_289),
	.R32(SYNTHESIZED_WIRE_290),
	.L1(SYNTHESIZED_WIRE_291),
	.L2(SYNTHESIZED_WIRE_292),
	.L3(SYNTHESIZED_WIRE_293),
	.L4(SYNTHESIZED_WIRE_294),
	.L5(SYNTHESIZED_WIRE_295),
	.L6(SYNTHESIZED_WIRE_296),
	.L7(SYNTHESIZED_WIRE_297),
	.L8(SYNTHESIZED_WIRE_298),
	.L9(SYNTHESIZED_WIRE_299),
	.L10(SYNTHESIZED_WIRE_300),
	.L11(SYNTHESIZED_WIRE_301),
	.L12(SYNTHESIZED_WIRE_302),
	.L13(SYNTHESIZED_WIRE_303),
	.L14(SYNTHESIZED_WIRE_304),
	.L15(SYNTHESIZED_WIRE_305),
	.L16(SYNTHESIZED_WIRE_306),
	.L17(SYNTHESIZED_WIRE_307),
	.L18(SYNTHESIZED_WIRE_308),
	.L19(SYNTHESIZED_WIRE_309),
	.L20(SYNTHESIZED_WIRE_310),
	.L21(SYNTHESIZED_WIRE_311),
	.L22(SYNTHESIZED_WIRE_312),
	.L23(SYNTHESIZED_WIRE_313),
	.L24(SYNTHESIZED_WIRE_314),
	.L25(SYNTHESIZED_WIRE_315),
	.L26(SYNTHESIZED_WIRE_316),
	.L27(SYNTHESIZED_WIRE_317),
	.L28(SYNTHESIZED_WIRE_318),
	.L29(SYNTHESIZED_WIRE_319),
	.L30(SYNTHESIZED_WIRE_320),
	.L31(SYNTHESIZED_WIRE_321),
	.L32(SYNTHESIZED_WIRE_322),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_323),
	.R_next1(SYNTHESIZED_WIRE_324),
	.R_next2(SYNTHESIZED_WIRE_325),
	.R_next3(SYNTHESIZED_WIRE_326),
	.R_next4(SYNTHESIZED_WIRE_327),
	.R_next5(SYNTHESIZED_WIRE_328),
	.R_next6(SYNTHESIZED_WIRE_329),
	.R_next7(SYNTHESIZED_WIRE_330),
	.R_next8(SYNTHESIZED_WIRE_331),
	.R_next9(SYNTHESIZED_WIRE_332),
	.R_next10(SYNTHESIZED_WIRE_333),
	.R_next11(SYNTHESIZED_WIRE_334),
	.R_next12(SYNTHESIZED_WIRE_335),
	.R_next13(SYNTHESIZED_WIRE_336),
	.R_next14(SYNTHESIZED_WIRE_337),
	.R_next15(SYNTHESIZED_WIRE_338),
	.R_next16(SYNTHESIZED_WIRE_339),
	.R_next17(SYNTHESIZED_WIRE_340),
	.R_next18(SYNTHESIZED_WIRE_341),
	.R_next19(SYNTHESIZED_WIRE_342),
	.R_next20(SYNTHESIZED_WIRE_343),
	.R_next21(SYNTHESIZED_WIRE_344),
	.R_next22(SYNTHESIZED_WIRE_345),
	.R_next23(SYNTHESIZED_WIRE_346),
	.R_next24(SYNTHESIZED_WIRE_347),
	.R_next25(SYNTHESIZED_WIRE_348),
	.R_next26(SYNTHESIZED_WIRE_349),
	.R_next27(SYNTHESIZED_WIRE_350),
	.R_next28(SYNTHESIZED_WIRE_351),
	.R_next29(SYNTHESIZED_WIRE_352),
	.R_next30(SYNTHESIZED_WIRE_353),
	.R_next31(SYNTHESIZED_WIRE_354),
	.R_next32(SYNTHESIZED_WIRE_355),
	.L_next1(SYNTHESIZED_WIRE_356),
	.L_next2(SYNTHESIZED_WIRE_357),
	.L_next3(SYNTHESIZED_WIRE_358),
	.L_next4(SYNTHESIZED_WIRE_359),
	.L_next5(SYNTHESIZED_WIRE_360),
	.L_next6(SYNTHESIZED_WIRE_361),
	.L_next7(SYNTHESIZED_WIRE_362),
	.L_next8(SYNTHESIZED_WIRE_363),
	.L_next9(SYNTHESIZED_WIRE_364),
	.L_next10(SYNTHESIZED_WIRE_365),
	.L_next11(SYNTHESIZED_WIRE_366),
	.L_next12(SYNTHESIZED_WIRE_367),
	.L_next13(SYNTHESIZED_WIRE_368),
	.L_next14(SYNTHESIZED_WIRE_369),
	.L_next15(SYNTHESIZED_WIRE_370),
	.L_next16(SYNTHESIZED_WIRE_371),
	.L_next17(SYNTHESIZED_WIRE_372),
	.L_next18(SYNTHESIZED_WIRE_373),
	.L_next19(SYNTHESIZED_WIRE_374),
	.L_next20(SYNTHESIZED_WIRE_375),
	.L_next21(SYNTHESIZED_WIRE_376),
	.L_next22(SYNTHESIZED_WIRE_377),
	.L_next23(SYNTHESIZED_WIRE_378),
	.L_next24(SYNTHESIZED_WIRE_379),
	.L_next25(SYNTHESIZED_WIRE_380),
	.L_next26(SYNTHESIZED_WIRE_381),
	.L_next27(SYNTHESIZED_WIRE_382),
	.L_next28(SYNTHESIZED_WIRE_383),
	.L_next29(SYNTHESIZED_WIRE_384),
	.L_next30(SYNTHESIZED_WIRE_385),
	.L_next31(SYNTHESIZED_WIRE_386),
	.L_next32(SYNTHESIZED_WIRE_387));


round	b2v_inst44(
	.R1(SYNTHESIZED_WIRE_324),
	.R2(SYNTHESIZED_WIRE_325),
	.R3(SYNTHESIZED_WIRE_326),
	.R4(SYNTHESIZED_WIRE_327),
	.R5(SYNTHESIZED_WIRE_328),
	.R6(SYNTHESIZED_WIRE_329),
	.R7(SYNTHESIZED_WIRE_330),
	.R8(SYNTHESIZED_WIRE_331),
	.R9(SYNTHESIZED_WIRE_332),
	.R10(SYNTHESIZED_WIRE_333),
	.R11(SYNTHESIZED_WIRE_334),
	.R12(SYNTHESIZED_WIRE_335),
	.R13(SYNTHESIZED_WIRE_336),
	.R14(SYNTHESIZED_WIRE_337),
	.R15(SYNTHESIZED_WIRE_338),
	.R16(SYNTHESIZED_WIRE_339),
	.R17(SYNTHESIZED_WIRE_340),
	.R18(SYNTHESIZED_WIRE_341),
	.R19(SYNTHESIZED_WIRE_342),
	.R20(SYNTHESIZED_WIRE_343),
	.R21(SYNTHESIZED_WIRE_344),
	.R22(SYNTHESIZED_WIRE_345),
	.R23(SYNTHESIZED_WIRE_346),
	.R24(SYNTHESIZED_WIRE_347),
	.R25(SYNTHESIZED_WIRE_348),
	.R26(SYNTHESIZED_WIRE_349),
	.R27(SYNTHESIZED_WIRE_350),
	.R28(SYNTHESIZED_WIRE_351),
	.R29(SYNTHESIZED_WIRE_352),
	.R30(SYNTHESIZED_WIRE_353),
	.R31(SYNTHESIZED_WIRE_354),
	.R32(SYNTHESIZED_WIRE_355),
	.L1(SYNTHESIZED_WIRE_356),
	.L2(SYNTHESIZED_WIRE_357),
	.L3(SYNTHESIZED_WIRE_358),
	.L4(SYNTHESIZED_WIRE_359),
	.L5(SYNTHESIZED_WIRE_360),
	.L6(SYNTHESIZED_WIRE_361),
	.L7(SYNTHESIZED_WIRE_362),
	.L8(SYNTHESIZED_WIRE_363),
	.L9(SYNTHESIZED_WIRE_364),
	.L10(SYNTHESIZED_WIRE_365),
	.L11(SYNTHESIZED_WIRE_366),
	.L12(SYNTHESIZED_WIRE_367),
	.L13(SYNTHESIZED_WIRE_368),
	.L14(SYNTHESIZED_WIRE_369),
	.L15(SYNTHESIZED_WIRE_370),
	.L16(SYNTHESIZED_WIRE_371),
	.L17(SYNTHESIZED_WIRE_372),
	.L18(SYNTHESIZED_WIRE_373),
	.L19(SYNTHESIZED_WIRE_374),
	.L20(SYNTHESIZED_WIRE_375),
	.L21(SYNTHESIZED_WIRE_376),
	.L22(SYNTHESIZED_WIRE_377),
	.L23(SYNTHESIZED_WIRE_378),
	.L24(SYNTHESIZED_WIRE_379),
	.L25(SYNTHESIZED_WIRE_380),
	.L26(SYNTHESIZED_WIRE_381),
	.L27(SYNTHESIZED_WIRE_382),
	.L28(SYNTHESIZED_WIRE_383),
	.L29(SYNTHESIZED_WIRE_384),
	.L30(SYNTHESIZED_WIRE_385),
	.L31(SYNTHESIZED_WIRE_386),
	.L32(SYNTHESIZED_WIRE_387),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_388),
	.R_next1(SYNTHESIZED_WIRE_389),
	.R_next2(SYNTHESIZED_WIRE_390),
	.R_next3(SYNTHESIZED_WIRE_391),
	.R_next4(SYNTHESIZED_WIRE_392),
	.R_next5(SYNTHESIZED_WIRE_393),
	.R_next6(SYNTHESIZED_WIRE_394),
	.R_next7(SYNTHESIZED_WIRE_395),
	.R_next8(SYNTHESIZED_WIRE_396),
	.R_next9(SYNTHESIZED_WIRE_397),
	.R_next10(SYNTHESIZED_WIRE_398),
	.R_next11(SYNTHESIZED_WIRE_399),
	.R_next12(SYNTHESIZED_WIRE_400),
	.R_next13(SYNTHESIZED_WIRE_401),
	.R_next14(SYNTHESIZED_WIRE_402),
	.R_next15(SYNTHESIZED_WIRE_403),
	.R_next16(SYNTHESIZED_WIRE_404),
	.R_next17(SYNTHESIZED_WIRE_405),
	.R_next18(SYNTHESIZED_WIRE_406),
	.R_next19(SYNTHESIZED_WIRE_407),
	.R_next20(SYNTHESIZED_WIRE_408),
	.R_next21(SYNTHESIZED_WIRE_409),
	.R_next22(SYNTHESIZED_WIRE_410),
	.R_next23(SYNTHESIZED_WIRE_411),
	.R_next24(SYNTHESIZED_WIRE_412),
	.R_next25(SYNTHESIZED_WIRE_413),
	.R_next26(SYNTHESIZED_WIRE_414),
	.R_next27(SYNTHESIZED_WIRE_415),
	.R_next28(SYNTHESIZED_WIRE_416),
	.R_next29(SYNTHESIZED_WIRE_417),
	.R_next30(SYNTHESIZED_WIRE_418),
	.R_next31(SYNTHESIZED_WIRE_419),
	.R_next32(SYNTHESIZED_WIRE_420),
	.L_next1(SYNTHESIZED_WIRE_421),
	.L_next2(SYNTHESIZED_WIRE_422),
	.L_next3(SYNTHESIZED_WIRE_423),
	.L_next4(SYNTHESIZED_WIRE_424),
	.L_next5(SYNTHESIZED_WIRE_425),
	.L_next6(SYNTHESIZED_WIRE_426),
	.L_next7(SYNTHESIZED_WIRE_427),
	.L_next8(SYNTHESIZED_WIRE_428),
	.L_next9(SYNTHESIZED_WIRE_429),
	.L_next10(SYNTHESIZED_WIRE_430),
	.L_next11(SYNTHESIZED_WIRE_431),
	.L_next12(SYNTHESIZED_WIRE_432),
	.L_next13(SYNTHESIZED_WIRE_433),
	.L_next14(SYNTHESIZED_WIRE_434),
	.L_next15(SYNTHESIZED_WIRE_435),
	.L_next16(SYNTHESIZED_WIRE_436),
	.L_next17(SYNTHESIZED_WIRE_437),
	.L_next18(SYNTHESIZED_WIRE_438),
	.L_next19(SYNTHESIZED_WIRE_439),
	.L_next20(SYNTHESIZED_WIRE_440),
	.L_next21(SYNTHESIZED_WIRE_441),
	.L_next22(SYNTHESIZED_WIRE_442),
	.L_next23(SYNTHESIZED_WIRE_443),
	.L_next24(SYNTHESIZED_WIRE_444),
	.L_next25(SYNTHESIZED_WIRE_445),
	.L_next26(SYNTHESIZED_WIRE_446),
	.L_next27(SYNTHESIZED_WIRE_447),
	.L_next28(SYNTHESIZED_WIRE_448),
	.L_next29(SYNTHESIZED_WIRE_449),
	.L_next30(SYNTHESIZED_WIRE_450),
	.L_next31(SYNTHESIZED_WIRE_451),
	.L_next32(SYNTHESIZED_WIRE_452));


round	b2v_inst45(
	.R1(SYNTHESIZED_WIRE_389),
	.R2(SYNTHESIZED_WIRE_390),
	.R3(SYNTHESIZED_WIRE_391),
	.R4(SYNTHESIZED_WIRE_392),
	.R5(SYNTHESIZED_WIRE_393),
	.R6(SYNTHESIZED_WIRE_394),
	.R7(SYNTHESIZED_WIRE_395),
	.R8(SYNTHESIZED_WIRE_396),
	.R9(SYNTHESIZED_WIRE_397),
	.R10(SYNTHESIZED_WIRE_398),
	.R11(SYNTHESIZED_WIRE_399),
	.R12(SYNTHESIZED_WIRE_400),
	.R13(SYNTHESIZED_WIRE_401),
	.R14(SYNTHESIZED_WIRE_402),
	.R15(SYNTHESIZED_WIRE_403),
	.R16(SYNTHESIZED_WIRE_404),
	.R17(SYNTHESIZED_WIRE_405),
	.R18(SYNTHESIZED_WIRE_406),
	.R19(SYNTHESIZED_WIRE_407),
	.R20(SYNTHESIZED_WIRE_408),
	.R21(SYNTHESIZED_WIRE_409),
	.R22(SYNTHESIZED_WIRE_410),
	.R23(SYNTHESIZED_WIRE_411),
	.R24(SYNTHESIZED_WIRE_412),
	.R25(SYNTHESIZED_WIRE_413),
	.R26(SYNTHESIZED_WIRE_414),
	.R27(SYNTHESIZED_WIRE_415),
	.R28(SYNTHESIZED_WIRE_416),
	.R29(SYNTHESIZED_WIRE_417),
	.R30(SYNTHESIZED_WIRE_418),
	.R31(SYNTHESIZED_WIRE_419),
	.R32(SYNTHESIZED_WIRE_420),
	.L1(SYNTHESIZED_WIRE_421),
	.L2(SYNTHESIZED_WIRE_422),
	.L3(SYNTHESIZED_WIRE_423),
	.L4(SYNTHESIZED_WIRE_424),
	.L5(SYNTHESIZED_WIRE_425),
	.L6(SYNTHESIZED_WIRE_426),
	.L7(SYNTHESIZED_WIRE_427),
	.L8(SYNTHESIZED_WIRE_428),
	.L9(SYNTHESIZED_WIRE_429),
	.L10(SYNTHESIZED_WIRE_430),
	.L11(SYNTHESIZED_WIRE_431),
	.L12(SYNTHESIZED_WIRE_432),
	.L13(SYNTHESIZED_WIRE_433),
	.L14(SYNTHESIZED_WIRE_434),
	.L15(SYNTHESIZED_WIRE_435),
	.L16(SYNTHESIZED_WIRE_436),
	.L17(SYNTHESIZED_WIRE_437),
	.L18(SYNTHESIZED_WIRE_438),
	.L19(SYNTHESIZED_WIRE_439),
	.L20(SYNTHESIZED_WIRE_440),
	.L21(SYNTHESIZED_WIRE_441),
	.L22(SYNTHESIZED_WIRE_442),
	.L23(SYNTHESIZED_WIRE_443),
	.L24(SYNTHESIZED_WIRE_444),
	.L25(SYNTHESIZED_WIRE_445),
	.L26(SYNTHESIZED_WIRE_446),
	.L27(SYNTHESIZED_WIRE_447),
	.L28(SYNTHESIZED_WIRE_448),
	.L29(SYNTHESIZED_WIRE_449),
	.L30(SYNTHESIZED_WIRE_450),
	.L31(SYNTHESIZED_WIRE_451),
	.L32(SYNTHESIZED_WIRE_452),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_453),
	.R_next1(SYNTHESIZED_WIRE_454),
	.R_next2(SYNTHESIZED_WIRE_455),
	.R_next3(SYNTHESIZED_WIRE_456),
	.R_next4(SYNTHESIZED_WIRE_457),
	.R_next5(SYNTHESIZED_WIRE_458),
	.R_next6(SYNTHESIZED_WIRE_459),
	.R_next7(SYNTHESIZED_WIRE_460),
	.R_next8(SYNTHESIZED_WIRE_461),
	.R_next9(SYNTHESIZED_WIRE_462),
	.R_next10(SYNTHESIZED_WIRE_463),
	.R_next11(SYNTHESIZED_WIRE_464),
	.R_next12(SYNTHESIZED_WIRE_465),
	.R_next13(SYNTHESIZED_WIRE_466),
	.R_next14(SYNTHESIZED_WIRE_467),
	.R_next15(SYNTHESIZED_WIRE_468),
	.R_next16(SYNTHESIZED_WIRE_469),
	.R_next17(SYNTHESIZED_WIRE_470),
	.R_next18(SYNTHESIZED_WIRE_471),
	.R_next19(SYNTHESIZED_WIRE_472),
	.R_next20(SYNTHESIZED_WIRE_473),
	.R_next21(SYNTHESIZED_WIRE_474),
	.R_next22(SYNTHESIZED_WIRE_475),
	.R_next23(SYNTHESIZED_WIRE_476),
	.R_next24(SYNTHESIZED_WIRE_477),
	.R_next25(SYNTHESIZED_WIRE_478),
	.R_next26(SYNTHESIZED_WIRE_479),
	.R_next27(SYNTHESIZED_WIRE_480),
	.R_next28(SYNTHESIZED_WIRE_481),
	.R_next29(SYNTHESIZED_WIRE_482),
	.R_next30(SYNTHESIZED_WIRE_483),
	.R_next31(SYNTHESIZED_WIRE_484),
	.R_next32(SYNTHESIZED_WIRE_485),
	.L_next1(SYNTHESIZED_WIRE_486),
	.L_next2(SYNTHESIZED_WIRE_487),
	.L_next3(SYNTHESIZED_WIRE_488),
	.L_next4(SYNTHESIZED_WIRE_489),
	.L_next5(SYNTHESIZED_WIRE_490),
	.L_next6(SYNTHESIZED_WIRE_491),
	.L_next7(SYNTHESIZED_WIRE_492),
	.L_next8(SYNTHESIZED_WIRE_493),
	.L_next9(SYNTHESIZED_WIRE_494),
	.L_next10(SYNTHESIZED_WIRE_495),
	.L_next11(SYNTHESIZED_WIRE_496),
	.L_next12(SYNTHESIZED_WIRE_497),
	.L_next13(SYNTHESIZED_WIRE_498),
	.L_next14(SYNTHESIZED_WIRE_499),
	.L_next15(SYNTHESIZED_WIRE_500),
	.L_next16(SYNTHESIZED_WIRE_501),
	.L_next17(SYNTHESIZED_WIRE_502),
	.L_next18(SYNTHESIZED_WIRE_503),
	.L_next19(SYNTHESIZED_WIRE_504),
	.L_next20(SYNTHESIZED_WIRE_505),
	.L_next21(SYNTHESIZED_WIRE_506),
	.L_next22(SYNTHESIZED_WIRE_507),
	.L_next23(SYNTHESIZED_WIRE_508),
	.L_next24(SYNTHESIZED_WIRE_509),
	.L_next25(SYNTHESIZED_WIRE_510),
	.L_next26(SYNTHESIZED_WIRE_511),
	.L_next27(SYNTHESIZED_WIRE_512),
	.L_next28(SYNTHESIZED_WIRE_513),
	.L_next29(SYNTHESIZED_WIRE_514),
	.L_next30(SYNTHESIZED_WIRE_515),
	.L_next31(SYNTHESIZED_WIRE_516),
	.L_next32(SYNTHESIZED_WIRE_517));


round	b2v_inst46(
	.R1(SYNTHESIZED_WIRE_454),
	.R2(SYNTHESIZED_WIRE_455),
	.R3(SYNTHESIZED_WIRE_456),
	.R4(SYNTHESIZED_WIRE_457),
	.R5(SYNTHESIZED_WIRE_458),
	.R6(SYNTHESIZED_WIRE_459),
	.R7(SYNTHESIZED_WIRE_460),
	.R8(SYNTHESIZED_WIRE_461),
	.R9(SYNTHESIZED_WIRE_462),
	.R10(SYNTHESIZED_WIRE_463),
	.R11(SYNTHESIZED_WIRE_464),
	.R12(SYNTHESIZED_WIRE_465),
	.R13(SYNTHESIZED_WIRE_466),
	.R14(SYNTHESIZED_WIRE_467),
	.R15(SYNTHESIZED_WIRE_468),
	.R16(SYNTHESIZED_WIRE_469),
	.R17(SYNTHESIZED_WIRE_470),
	.R18(SYNTHESIZED_WIRE_471),
	.R19(SYNTHESIZED_WIRE_472),
	.R20(SYNTHESIZED_WIRE_473),
	.R21(SYNTHESIZED_WIRE_474),
	.R22(SYNTHESIZED_WIRE_475),
	.R23(SYNTHESIZED_WIRE_476),
	.R24(SYNTHESIZED_WIRE_477),
	.R25(SYNTHESIZED_WIRE_478),
	.R26(SYNTHESIZED_WIRE_479),
	.R27(SYNTHESIZED_WIRE_480),
	.R28(SYNTHESIZED_WIRE_481),
	.R29(SYNTHESIZED_WIRE_482),
	.R30(SYNTHESIZED_WIRE_483),
	.R31(SYNTHESIZED_WIRE_484),
	.R32(SYNTHESIZED_WIRE_485),
	.L1(SYNTHESIZED_WIRE_486),
	.L2(SYNTHESIZED_WIRE_487),
	.L3(SYNTHESIZED_WIRE_488),
	.L4(SYNTHESIZED_WIRE_489),
	.L5(SYNTHESIZED_WIRE_490),
	.L6(SYNTHESIZED_WIRE_491),
	.L7(SYNTHESIZED_WIRE_492),
	.L8(SYNTHESIZED_WIRE_493),
	.L9(SYNTHESIZED_WIRE_494),
	.L10(SYNTHESIZED_WIRE_495),
	.L11(SYNTHESIZED_WIRE_496),
	.L12(SYNTHESIZED_WIRE_497),
	.L13(SYNTHESIZED_WIRE_498),
	.L14(SYNTHESIZED_WIRE_499),
	.L15(SYNTHESIZED_WIRE_500),
	.L16(SYNTHESIZED_WIRE_501),
	.L17(SYNTHESIZED_WIRE_502),
	.L18(SYNTHESIZED_WIRE_503),
	.L19(SYNTHESIZED_WIRE_504),
	.L20(SYNTHESIZED_WIRE_505),
	.L21(SYNTHESIZED_WIRE_506),
	.L22(SYNTHESIZED_WIRE_507),
	.L23(SYNTHESIZED_WIRE_508),
	.L24(SYNTHESIZED_WIRE_509),
	.L25(SYNTHESIZED_WIRE_510),
	.L26(SYNTHESIZED_WIRE_511),
	.L27(SYNTHESIZED_WIRE_512),
	.L28(SYNTHESIZED_WIRE_513),
	.L29(SYNTHESIZED_WIRE_514),
	.L30(SYNTHESIZED_WIRE_515),
	.L31(SYNTHESIZED_WIRE_516),
	.L32(SYNTHESIZED_WIRE_517),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_518),
	.R_next1(SYNTHESIZED_WIRE_519),
	.R_next2(SYNTHESIZED_WIRE_520),
	.R_next3(SYNTHESIZED_WIRE_521),
	.R_next4(SYNTHESIZED_WIRE_522),
	.R_next5(SYNTHESIZED_WIRE_523),
	.R_next6(SYNTHESIZED_WIRE_524),
	.R_next7(SYNTHESIZED_WIRE_525),
	.R_next8(SYNTHESIZED_WIRE_526),
	.R_next9(SYNTHESIZED_WIRE_527),
	.R_next10(SYNTHESIZED_WIRE_528),
	.R_next11(SYNTHESIZED_WIRE_529),
	.R_next12(SYNTHESIZED_WIRE_530),
	.R_next13(SYNTHESIZED_WIRE_531),
	.R_next14(SYNTHESIZED_WIRE_532),
	.R_next15(SYNTHESIZED_WIRE_533),
	.R_next16(SYNTHESIZED_WIRE_534),
	.R_next17(SYNTHESIZED_WIRE_535),
	.R_next18(SYNTHESIZED_WIRE_536),
	.R_next19(SYNTHESIZED_WIRE_537),
	.R_next20(SYNTHESIZED_WIRE_538),
	.R_next21(SYNTHESIZED_WIRE_539),
	.R_next22(SYNTHESIZED_WIRE_540),
	.R_next23(SYNTHESIZED_WIRE_541),
	.R_next24(SYNTHESIZED_WIRE_542),
	.R_next25(SYNTHESIZED_WIRE_543),
	.R_next26(SYNTHESIZED_WIRE_544),
	.R_next27(SYNTHESIZED_WIRE_545),
	.R_next28(SYNTHESIZED_WIRE_546),
	.R_next29(SYNTHESIZED_WIRE_547),
	.R_next30(SYNTHESIZED_WIRE_548),
	.R_next31(SYNTHESIZED_WIRE_549),
	.R_next32(SYNTHESIZED_WIRE_550),
	.L_next1(SYNTHESIZED_WIRE_551),
	.L_next2(SYNTHESIZED_WIRE_552),
	.L_next3(SYNTHESIZED_WIRE_553),
	.L_next4(SYNTHESIZED_WIRE_554),
	.L_next5(SYNTHESIZED_WIRE_555),
	.L_next6(SYNTHESIZED_WIRE_556),
	.L_next7(SYNTHESIZED_WIRE_557),
	.L_next8(SYNTHESIZED_WIRE_558),
	.L_next9(SYNTHESIZED_WIRE_559),
	.L_next10(SYNTHESIZED_WIRE_560),
	.L_next11(SYNTHESIZED_WIRE_561),
	.L_next12(SYNTHESIZED_WIRE_562),
	.L_next13(SYNTHESIZED_WIRE_563),
	.L_next14(SYNTHESIZED_WIRE_564),
	.L_next15(SYNTHESIZED_WIRE_565),
	.L_next16(SYNTHESIZED_WIRE_566),
	.L_next17(SYNTHESIZED_WIRE_567),
	.L_next18(SYNTHESIZED_WIRE_568),
	.L_next19(SYNTHESIZED_WIRE_569),
	.L_next20(SYNTHESIZED_WIRE_570),
	.L_next21(SYNTHESIZED_WIRE_571),
	.L_next22(SYNTHESIZED_WIRE_572),
	.L_next23(SYNTHESIZED_WIRE_573),
	.L_next24(SYNTHESIZED_WIRE_574),
	.L_next25(SYNTHESIZED_WIRE_575),
	.L_next26(SYNTHESIZED_WIRE_576),
	.L_next27(SYNTHESIZED_WIRE_577),
	.L_next28(SYNTHESIZED_WIRE_578),
	.L_next29(SYNTHESIZED_WIRE_579),
	.L_next30(SYNTHESIZED_WIRE_580),
	.L_next31(SYNTHESIZED_WIRE_581),
	.L_next32(SYNTHESIZED_WIRE_582));


round	b2v_inst47(
	.R1(SYNTHESIZED_WIRE_519),
	.R2(SYNTHESIZED_WIRE_520),
	.R3(SYNTHESIZED_WIRE_521),
	.R4(SYNTHESIZED_WIRE_522),
	.R5(SYNTHESIZED_WIRE_523),
	.R6(SYNTHESIZED_WIRE_524),
	.R7(SYNTHESIZED_WIRE_525),
	.R8(SYNTHESIZED_WIRE_526),
	.R9(SYNTHESIZED_WIRE_527),
	.R10(SYNTHESIZED_WIRE_528),
	.R11(SYNTHESIZED_WIRE_529),
	.R12(SYNTHESIZED_WIRE_530),
	.R13(SYNTHESIZED_WIRE_531),
	.R14(SYNTHESIZED_WIRE_532),
	.R15(SYNTHESIZED_WIRE_533),
	.R16(SYNTHESIZED_WIRE_534),
	.R17(SYNTHESIZED_WIRE_535),
	.R18(SYNTHESIZED_WIRE_536),
	.R19(SYNTHESIZED_WIRE_537),
	.R20(SYNTHESIZED_WIRE_538),
	.R21(SYNTHESIZED_WIRE_539),
	.R22(SYNTHESIZED_WIRE_540),
	.R23(SYNTHESIZED_WIRE_541),
	.R24(SYNTHESIZED_WIRE_542),
	.R25(SYNTHESIZED_WIRE_543),
	.R26(SYNTHESIZED_WIRE_544),
	.R27(SYNTHESIZED_WIRE_545),
	.R28(SYNTHESIZED_WIRE_546),
	.R29(SYNTHESIZED_WIRE_547),
	.R30(SYNTHESIZED_WIRE_548),
	.R31(SYNTHESIZED_WIRE_549),
	.R32(SYNTHESIZED_WIRE_550),
	.L1(SYNTHESIZED_WIRE_551),
	.L2(SYNTHESIZED_WIRE_552),
	.L3(SYNTHESIZED_WIRE_553),
	.L4(SYNTHESIZED_WIRE_554),
	.L5(SYNTHESIZED_WIRE_555),
	.L6(SYNTHESIZED_WIRE_556),
	.L7(SYNTHESIZED_WIRE_557),
	.L8(SYNTHESIZED_WIRE_558),
	.L9(SYNTHESIZED_WIRE_559),
	.L10(SYNTHESIZED_WIRE_560),
	.L11(SYNTHESIZED_WIRE_561),
	.L12(SYNTHESIZED_WIRE_562),
	.L13(SYNTHESIZED_WIRE_563),
	.L14(SYNTHESIZED_WIRE_564),
	.L15(SYNTHESIZED_WIRE_565),
	.L16(SYNTHESIZED_WIRE_566),
	.L17(SYNTHESIZED_WIRE_567),
	.L18(SYNTHESIZED_WIRE_568),
	.L19(SYNTHESIZED_WIRE_569),
	.L20(SYNTHESIZED_WIRE_570),
	.L21(SYNTHESIZED_WIRE_571),
	.L22(SYNTHESIZED_WIRE_572),
	.L23(SYNTHESIZED_WIRE_573),
	.L24(SYNTHESIZED_WIRE_574),
	.L25(SYNTHESIZED_WIRE_575),
	.L26(SYNTHESIZED_WIRE_576),
	.L27(SYNTHESIZED_WIRE_577),
	.L28(SYNTHESIZED_WIRE_578),
	.L29(SYNTHESIZED_WIRE_579),
	.L30(SYNTHESIZED_WIRE_580),
	.L31(SYNTHESIZED_WIRE_581),
	.L32(SYNTHESIZED_WIRE_582),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_583),
	.R_next1(SYNTHESIZED_WIRE_584),
	.R_next2(SYNTHESIZED_WIRE_585),
	.R_next3(SYNTHESIZED_WIRE_586),
	.R_next4(SYNTHESIZED_WIRE_587),
	.R_next5(SYNTHESIZED_WIRE_588),
	.R_next6(SYNTHESIZED_WIRE_589),
	.R_next7(SYNTHESIZED_WIRE_590),
	.R_next8(SYNTHESIZED_WIRE_591),
	.R_next9(SYNTHESIZED_WIRE_592),
	.R_next10(SYNTHESIZED_WIRE_593),
	.R_next11(SYNTHESIZED_WIRE_594),
	.R_next12(SYNTHESIZED_WIRE_595),
	.R_next13(SYNTHESIZED_WIRE_596),
	.R_next14(SYNTHESIZED_WIRE_597),
	.R_next15(SYNTHESIZED_WIRE_598),
	.R_next16(SYNTHESIZED_WIRE_599),
	.R_next17(SYNTHESIZED_WIRE_600),
	.R_next18(SYNTHESIZED_WIRE_601),
	.R_next19(SYNTHESIZED_WIRE_602),
	.R_next20(SYNTHESIZED_WIRE_603),
	.R_next21(SYNTHESIZED_WIRE_604),
	.R_next22(SYNTHESIZED_WIRE_605),
	.R_next23(SYNTHESIZED_WIRE_606),
	.R_next24(SYNTHESIZED_WIRE_607),
	.R_next25(SYNTHESIZED_WIRE_608),
	.R_next26(SYNTHESIZED_WIRE_609),
	.R_next27(SYNTHESIZED_WIRE_610),
	.R_next28(SYNTHESIZED_WIRE_611),
	.R_next29(SYNTHESIZED_WIRE_612),
	.R_next30(SYNTHESIZED_WIRE_613),
	.R_next31(SYNTHESIZED_WIRE_614),
	.R_next32(SYNTHESIZED_WIRE_615),
	.L_next1(SYNTHESIZED_WIRE_616),
	.L_next2(SYNTHESIZED_WIRE_617),
	.L_next3(SYNTHESIZED_WIRE_618),
	.L_next4(SYNTHESIZED_WIRE_619),
	.L_next5(SYNTHESIZED_WIRE_620),
	.L_next6(SYNTHESIZED_WIRE_621),
	.L_next7(SYNTHESIZED_WIRE_622),
	.L_next8(SYNTHESIZED_WIRE_623),
	.L_next9(SYNTHESIZED_WIRE_624),
	.L_next10(SYNTHESIZED_WIRE_625),
	.L_next11(SYNTHESIZED_WIRE_626),
	.L_next12(SYNTHESIZED_WIRE_627),
	.L_next13(SYNTHESIZED_WIRE_628),
	.L_next14(SYNTHESIZED_WIRE_629),
	.L_next15(SYNTHESIZED_WIRE_630),
	.L_next16(SYNTHESIZED_WIRE_631),
	.L_next17(SYNTHESIZED_WIRE_632),
	.L_next18(SYNTHESIZED_WIRE_633),
	.L_next19(SYNTHESIZED_WIRE_634),
	.L_next20(SYNTHESIZED_WIRE_635),
	.L_next21(SYNTHESIZED_WIRE_636),
	.L_next22(SYNTHESIZED_WIRE_637),
	.L_next23(SYNTHESIZED_WIRE_638),
	.L_next24(SYNTHESIZED_WIRE_639),
	.L_next25(SYNTHESIZED_WIRE_640),
	.L_next26(SYNTHESIZED_WIRE_641),
	.L_next27(SYNTHESIZED_WIRE_642),
	.L_next28(SYNTHESIZED_WIRE_643),
	.L_next29(SYNTHESIZED_WIRE_644),
	.L_next30(SYNTHESIZED_WIRE_645),
	.L_next31(SYNTHESIZED_WIRE_646),
	.L_next32(SYNTHESIZED_WIRE_647));


round	b2v_inst48(
	.R1(SYNTHESIZED_WIRE_584),
	.R2(SYNTHESIZED_WIRE_585),
	.R3(SYNTHESIZED_WIRE_586),
	.R4(SYNTHESIZED_WIRE_587),
	.R5(SYNTHESIZED_WIRE_588),
	.R6(SYNTHESIZED_WIRE_589),
	.R7(SYNTHESIZED_WIRE_590),
	.R8(SYNTHESIZED_WIRE_591),
	.R9(SYNTHESIZED_WIRE_592),
	.R10(SYNTHESIZED_WIRE_593),
	.R11(SYNTHESIZED_WIRE_594),
	.R12(SYNTHESIZED_WIRE_595),
	.R13(SYNTHESIZED_WIRE_596),
	.R14(SYNTHESIZED_WIRE_597),
	.R15(SYNTHESIZED_WIRE_598),
	.R16(SYNTHESIZED_WIRE_599),
	.R17(SYNTHESIZED_WIRE_600),
	.R18(SYNTHESIZED_WIRE_601),
	.R19(SYNTHESIZED_WIRE_602),
	.R20(SYNTHESIZED_WIRE_603),
	.R21(SYNTHESIZED_WIRE_604),
	.R22(SYNTHESIZED_WIRE_605),
	.R23(SYNTHESIZED_WIRE_606),
	.R24(SYNTHESIZED_WIRE_607),
	.R25(SYNTHESIZED_WIRE_608),
	.R26(SYNTHESIZED_WIRE_609),
	.R27(SYNTHESIZED_WIRE_610),
	.R28(SYNTHESIZED_WIRE_611),
	.R29(SYNTHESIZED_WIRE_612),
	.R30(SYNTHESIZED_WIRE_613),
	.R31(SYNTHESIZED_WIRE_614),
	.R32(SYNTHESIZED_WIRE_615),
	.L1(SYNTHESIZED_WIRE_616),
	.L2(SYNTHESIZED_WIRE_617),
	.L3(SYNTHESIZED_WIRE_618),
	.L4(SYNTHESIZED_WIRE_619),
	.L5(SYNTHESIZED_WIRE_620),
	.L6(SYNTHESIZED_WIRE_621),
	.L7(SYNTHESIZED_WIRE_622),
	.L8(SYNTHESIZED_WIRE_623),
	.L9(SYNTHESIZED_WIRE_624),
	.L10(SYNTHESIZED_WIRE_625),
	.L11(SYNTHESIZED_WIRE_626),
	.L12(SYNTHESIZED_WIRE_627),
	.L13(SYNTHESIZED_WIRE_628),
	.L14(SYNTHESIZED_WIRE_629),
	.L15(SYNTHESIZED_WIRE_630),
	.L16(SYNTHESIZED_WIRE_631),
	.L17(SYNTHESIZED_WIRE_632),
	.L18(SYNTHESIZED_WIRE_633),
	.L19(SYNTHESIZED_WIRE_634),
	.L20(SYNTHESIZED_WIRE_635),
	.L21(SYNTHESIZED_WIRE_636),
	.L22(SYNTHESIZED_WIRE_637),
	.L23(SYNTHESIZED_WIRE_638),
	.L24(SYNTHESIZED_WIRE_639),
	.L25(SYNTHESIZED_WIRE_640),
	.L26(SYNTHESIZED_WIRE_641),
	.L27(SYNTHESIZED_WIRE_642),
	.L28(SYNTHESIZED_WIRE_643),
	.L29(SYNTHESIZED_WIRE_644),
	.L30(SYNTHESIZED_WIRE_645),
	.L31(SYNTHESIZED_WIRE_646),
	.L32(SYNTHESIZED_WIRE_647),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_648),
	.R_next1(SYNTHESIZED_WIRE_649),
	.R_next2(SYNTHESIZED_WIRE_650),
	.R_next3(SYNTHESIZED_WIRE_651),
	.R_next4(SYNTHESIZED_WIRE_652),
	.R_next5(SYNTHESIZED_WIRE_653),
	.R_next6(SYNTHESIZED_WIRE_654),
	.R_next7(SYNTHESIZED_WIRE_655),
	.R_next8(SYNTHESIZED_WIRE_656),
	.R_next9(SYNTHESIZED_WIRE_657),
	.R_next10(SYNTHESIZED_WIRE_658),
	.R_next11(SYNTHESIZED_WIRE_659),
	.R_next12(SYNTHESIZED_WIRE_660),
	.R_next13(SYNTHESIZED_WIRE_661),
	.R_next14(SYNTHESIZED_WIRE_662),
	.R_next15(SYNTHESIZED_WIRE_663),
	.R_next16(SYNTHESIZED_WIRE_664),
	.R_next17(SYNTHESIZED_WIRE_665),
	.R_next18(SYNTHESIZED_WIRE_666),
	.R_next19(SYNTHESIZED_WIRE_667),
	.R_next20(SYNTHESIZED_WIRE_668),
	.R_next21(SYNTHESIZED_WIRE_669),
	.R_next22(SYNTHESIZED_WIRE_670),
	.R_next23(SYNTHESIZED_WIRE_671),
	.R_next24(SYNTHESIZED_WIRE_672),
	.R_next25(SYNTHESIZED_WIRE_673),
	.R_next26(SYNTHESIZED_WIRE_674),
	.R_next27(SYNTHESIZED_WIRE_675),
	.R_next28(SYNTHESIZED_WIRE_676),
	.R_next29(SYNTHESIZED_WIRE_677),
	.R_next30(SYNTHESIZED_WIRE_678),
	.R_next31(SYNTHESIZED_WIRE_679),
	.R_next32(SYNTHESIZED_WIRE_680),
	.L_next1(SYNTHESIZED_WIRE_681),
	.L_next2(SYNTHESIZED_WIRE_682),
	.L_next3(SYNTHESIZED_WIRE_683),
	.L_next4(SYNTHESIZED_WIRE_684),
	.L_next5(SYNTHESIZED_WIRE_685),
	.L_next6(SYNTHESIZED_WIRE_686),
	.L_next7(SYNTHESIZED_WIRE_687),
	.L_next8(SYNTHESIZED_WIRE_688),
	.L_next9(SYNTHESIZED_WIRE_689),
	.L_next10(SYNTHESIZED_WIRE_690),
	.L_next11(SYNTHESIZED_WIRE_691),
	.L_next12(SYNTHESIZED_WIRE_692),
	.L_next13(SYNTHESIZED_WIRE_693),
	.L_next14(SYNTHESIZED_WIRE_694),
	.L_next15(SYNTHESIZED_WIRE_695),
	.L_next16(SYNTHESIZED_WIRE_696),
	.L_next17(SYNTHESIZED_WIRE_697),
	.L_next18(SYNTHESIZED_WIRE_698),
	.L_next19(SYNTHESIZED_WIRE_699),
	.L_next20(SYNTHESIZED_WIRE_700),
	.L_next21(SYNTHESIZED_WIRE_701),
	.L_next22(SYNTHESIZED_WIRE_702),
	.L_next23(SYNTHESIZED_WIRE_703),
	.L_next24(SYNTHESIZED_WIRE_704),
	.L_next25(SYNTHESIZED_WIRE_705),
	.L_next26(SYNTHESIZED_WIRE_706),
	.L_next27(SYNTHESIZED_WIRE_707),
	.L_next28(SYNTHESIZED_WIRE_708),
	.L_next29(SYNTHESIZED_WIRE_709),
	.L_next30(SYNTHESIZED_WIRE_710),
	.L_next31(SYNTHESIZED_WIRE_711),
	.L_next32(SYNTHESIZED_WIRE_712));


round	b2v_inst49(
	.R1(SYNTHESIZED_WIRE_649),
	.R2(SYNTHESIZED_WIRE_650),
	.R3(SYNTHESIZED_WIRE_651),
	.R4(SYNTHESIZED_WIRE_652),
	.R5(SYNTHESIZED_WIRE_653),
	.R6(SYNTHESIZED_WIRE_654),
	.R7(SYNTHESIZED_WIRE_655),
	.R8(SYNTHESIZED_WIRE_656),
	.R9(SYNTHESIZED_WIRE_657),
	.R10(SYNTHESIZED_WIRE_658),
	.R11(SYNTHESIZED_WIRE_659),
	.R12(SYNTHESIZED_WIRE_660),
	.R13(SYNTHESIZED_WIRE_661),
	.R14(SYNTHESIZED_WIRE_662),
	.R15(SYNTHESIZED_WIRE_663),
	.R16(SYNTHESIZED_WIRE_664),
	.R17(SYNTHESIZED_WIRE_665),
	.R18(SYNTHESIZED_WIRE_666),
	.R19(SYNTHESIZED_WIRE_667),
	.R20(SYNTHESIZED_WIRE_668),
	.R21(SYNTHESIZED_WIRE_669),
	.R22(SYNTHESIZED_WIRE_670),
	.R23(SYNTHESIZED_WIRE_671),
	.R24(SYNTHESIZED_WIRE_672),
	.R25(SYNTHESIZED_WIRE_673),
	.R26(SYNTHESIZED_WIRE_674),
	.R27(SYNTHESIZED_WIRE_675),
	.R28(SYNTHESIZED_WIRE_676),
	.R29(SYNTHESIZED_WIRE_677),
	.R30(SYNTHESIZED_WIRE_678),
	.R31(SYNTHESIZED_WIRE_679),
	.R32(SYNTHESIZED_WIRE_680),
	.L1(SYNTHESIZED_WIRE_681),
	.L2(SYNTHESIZED_WIRE_682),
	.L3(SYNTHESIZED_WIRE_683),
	.L4(SYNTHESIZED_WIRE_684),
	.L5(SYNTHESIZED_WIRE_685),
	.L6(SYNTHESIZED_WIRE_686),
	.L7(SYNTHESIZED_WIRE_687),
	.L8(SYNTHESIZED_WIRE_688),
	.L9(SYNTHESIZED_WIRE_689),
	.L10(SYNTHESIZED_WIRE_690),
	.L11(SYNTHESIZED_WIRE_691),
	.L12(SYNTHESIZED_WIRE_692),
	.L13(SYNTHESIZED_WIRE_693),
	.L14(SYNTHESIZED_WIRE_694),
	.L15(SYNTHESIZED_WIRE_695),
	.L16(SYNTHESIZED_WIRE_696),
	.L17(SYNTHESIZED_WIRE_697),
	.L18(SYNTHESIZED_WIRE_698),
	.L19(SYNTHESIZED_WIRE_699),
	.L20(SYNTHESIZED_WIRE_700),
	.L21(SYNTHESIZED_WIRE_701),
	.L22(SYNTHESIZED_WIRE_702),
	.L23(SYNTHESIZED_WIRE_703),
	.L24(SYNTHESIZED_WIRE_704),
	.L25(SYNTHESIZED_WIRE_705),
	.L26(SYNTHESIZED_WIRE_706),
	.L27(SYNTHESIZED_WIRE_707),
	.L28(SYNTHESIZED_WIRE_708),
	.L29(SYNTHESIZED_WIRE_709),
	.L30(SYNTHESIZED_WIRE_710),
	.L31(SYNTHESIZED_WIRE_711),
	.L32(SYNTHESIZED_WIRE_712),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_713),
	.R_next1(SYNTHESIZED_WIRE_714),
	.R_next2(SYNTHESIZED_WIRE_715),
	.R_next3(SYNTHESIZED_WIRE_716),
	.R_next4(SYNTHESIZED_WIRE_717),
	.R_next5(SYNTHESIZED_WIRE_718),
	.R_next6(SYNTHESIZED_WIRE_719),
	.R_next7(SYNTHESIZED_WIRE_720),
	.R_next8(SYNTHESIZED_WIRE_721),
	.R_next9(SYNTHESIZED_WIRE_722),
	.R_next10(SYNTHESIZED_WIRE_723),
	.R_next11(SYNTHESIZED_WIRE_724),
	.R_next12(SYNTHESIZED_WIRE_725),
	.R_next13(SYNTHESIZED_WIRE_726),
	.R_next14(SYNTHESIZED_WIRE_727),
	.R_next15(SYNTHESIZED_WIRE_728),
	.R_next16(SYNTHESIZED_WIRE_729),
	.R_next17(SYNTHESIZED_WIRE_730),
	.R_next18(SYNTHESIZED_WIRE_731),
	.R_next19(SYNTHESIZED_WIRE_732),
	.R_next20(SYNTHESIZED_WIRE_733),
	.R_next21(SYNTHESIZED_WIRE_734),
	.R_next22(SYNTHESIZED_WIRE_735),
	.R_next23(SYNTHESIZED_WIRE_736),
	.R_next24(SYNTHESIZED_WIRE_737),
	.R_next25(SYNTHESIZED_WIRE_738),
	.R_next26(SYNTHESIZED_WIRE_739),
	.R_next27(SYNTHESIZED_WIRE_740),
	.R_next28(SYNTHESIZED_WIRE_741),
	.R_next29(SYNTHESIZED_WIRE_742),
	.R_next30(SYNTHESIZED_WIRE_743),
	.R_next31(SYNTHESIZED_WIRE_744),
	.R_next32(SYNTHESIZED_WIRE_745),
	.L_next1(SYNTHESIZED_WIRE_746),
	.L_next2(SYNTHESIZED_WIRE_747),
	.L_next3(SYNTHESIZED_WIRE_748),
	.L_next4(SYNTHESIZED_WIRE_749),
	.L_next5(SYNTHESIZED_WIRE_750),
	.L_next6(SYNTHESIZED_WIRE_751),
	.L_next7(SYNTHESIZED_WIRE_752),
	.L_next8(SYNTHESIZED_WIRE_753),
	.L_next9(SYNTHESIZED_WIRE_754),
	.L_next10(SYNTHESIZED_WIRE_755),
	.L_next11(SYNTHESIZED_WIRE_756),
	.L_next12(SYNTHESIZED_WIRE_757),
	.L_next13(SYNTHESIZED_WIRE_758),
	.L_next14(SYNTHESIZED_WIRE_759),
	.L_next15(SYNTHESIZED_WIRE_760),
	.L_next16(SYNTHESIZED_WIRE_761),
	.L_next17(SYNTHESIZED_WIRE_762),
	.L_next18(SYNTHESIZED_WIRE_763),
	.L_next19(SYNTHESIZED_WIRE_764),
	.L_next20(SYNTHESIZED_WIRE_765),
	.L_next21(SYNTHESIZED_WIRE_766),
	.L_next22(SYNTHESIZED_WIRE_767),
	.L_next23(SYNTHESIZED_WIRE_768),
	.L_next24(SYNTHESIZED_WIRE_769),
	.L_next25(SYNTHESIZED_WIRE_770),
	.L_next26(SYNTHESIZED_WIRE_771),
	.L_next27(SYNTHESIZED_WIRE_772),
	.L_next28(SYNTHESIZED_WIRE_773),
	.L_next29(SYNTHESIZED_WIRE_774),
	.L_next30(SYNTHESIZED_WIRE_775),
	.L_next31(SYNTHESIZED_WIRE_776),
	.L_next32(SYNTHESIZED_WIRE_777));


round	b2v_inst50(
	.R1(SYNTHESIZED_WIRE_714),
	.R2(SYNTHESIZED_WIRE_715),
	.R3(SYNTHESIZED_WIRE_716),
	.R4(SYNTHESIZED_WIRE_717),
	.R5(SYNTHESIZED_WIRE_718),
	.R6(SYNTHESIZED_WIRE_719),
	.R7(SYNTHESIZED_WIRE_720),
	.R8(SYNTHESIZED_WIRE_721),
	.R9(SYNTHESIZED_WIRE_722),
	.R10(SYNTHESIZED_WIRE_723),
	.R11(SYNTHESIZED_WIRE_724),
	.R12(SYNTHESIZED_WIRE_725),
	.R13(SYNTHESIZED_WIRE_726),
	.R14(SYNTHESIZED_WIRE_727),
	.R15(SYNTHESIZED_WIRE_728),
	.R16(SYNTHESIZED_WIRE_729),
	.R17(SYNTHESIZED_WIRE_730),
	.R18(SYNTHESIZED_WIRE_731),
	.R19(SYNTHESIZED_WIRE_732),
	.R20(SYNTHESIZED_WIRE_733),
	.R21(SYNTHESIZED_WIRE_734),
	.R22(SYNTHESIZED_WIRE_735),
	.R23(SYNTHESIZED_WIRE_736),
	.R24(SYNTHESIZED_WIRE_737),
	.R25(SYNTHESIZED_WIRE_738),
	.R26(SYNTHESIZED_WIRE_739),
	.R27(SYNTHESIZED_WIRE_740),
	.R28(SYNTHESIZED_WIRE_741),
	.R29(SYNTHESIZED_WIRE_742),
	.R30(SYNTHESIZED_WIRE_743),
	.R31(SYNTHESIZED_WIRE_744),
	.R32(SYNTHESIZED_WIRE_745),
	.L1(SYNTHESIZED_WIRE_746),
	.L2(SYNTHESIZED_WIRE_747),
	.L3(SYNTHESIZED_WIRE_748),
	.L4(SYNTHESIZED_WIRE_749),
	.L5(SYNTHESIZED_WIRE_750),
	.L6(SYNTHESIZED_WIRE_751),
	.L7(SYNTHESIZED_WIRE_752),
	.L8(SYNTHESIZED_WIRE_753),
	.L9(SYNTHESIZED_WIRE_754),
	.L10(SYNTHESIZED_WIRE_755),
	.L11(SYNTHESIZED_WIRE_756),
	.L12(SYNTHESIZED_WIRE_757),
	.L13(SYNTHESIZED_WIRE_758),
	.L14(SYNTHESIZED_WIRE_759),
	.L15(SYNTHESIZED_WIRE_760),
	.L16(SYNTHESIZED_WIRE_761),
	.L17(SYNTHESIZED_WIRE_762),
	.L18(SYNTHESIZED_WIRE_763),
	.L19(SYNTHESIZED_WIRE_764),
	.L20(SYNTHESIZED_WIRE_765),
	.L21(SYNTHESIZED_WIRE_766),
	.L22(SYNTHESIZED_WIRE_767),
	.L23(SYNTHESIZED_WIRE_768),
	.L24(SYNTHESIZED_WIRE_769),
	.L25(SYNTHESIZED_WIRE_770),
	.L26(SYNTHESIZED_WIRE_771),
	.L27(SYNTHESIZED_WIRE_772),
	.L28(SYNTHESIZED_WIRE_773),
	.L29(SYNTHESIZED_WIRE_774),
	.L30(SYNTHESIZED_WIRE_775),
	.L31(SYNTHESIZED_WIRE_776),
	.L32(SYNTHESIZED_WIRE_777),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_778),
	.R_next1(SYNTHESIZED_WIRE_779),
	.R_next2(SYNTHESIZED_WIRE_780),
	.R_next3(SYNTHESIZED_WIRE_781),
	.R_next4(SYNTHESIZED_WIRE_782),
	.R_next5(SYNTHESIZED_WIRE_783),
	.R_next6(SYNTHESIZED_WIRE_784),
	.R_next7(SYNTHESIZED_WIRE_785),
	.R_next8(SYNTHESIZED_WIRE_786),
	.R_next9(SYNTHESIZED_WIRE_787),
	.R_next10(SYNTHESIZED_WIRE_788),
	.R_next11(SYNTHESIZED_WIRE_789),
	.R_next12(SYNTHESIZED_WIRE_790),
	.R_next13(SYNTHESIZED_WIRE_791),
	.R_next14(SYNTHESIZED_WIRE_792),
	.R_next15(SYNTHESIZED_WIRE_793),
	.R_next16(SYNTHESIZED_WIRE_794),
	.R_next17(SYNTHESIZED_WIRE_795),
	.R_next18(SYNTHESIZED_WIRE_796),
	.R_next19(SYNTHESIZED_WIRE_797),
	.R_next20(SYNTHESIZED_WIRE_798),
	.R_next21(SYNTHESIZED_WIRE_799),
	.R_next22(SYNTHESIZED_WIRE_800),
	.R_next23(SYNTHESIZED_WIRE_801),
	.R_next24(SYNTHESIZED_WIRE_802),
	.R_next25(SYNTHESIZED_WIRE_803),
	.R_next26(SYNTHESIZED_WIRE_804),
	.R_next27(SYNTHESIZED_WIRE_805),
	.R_next28(SYNTHESIZED_WIRE_806),
	.R_next29(SYNTHESIZED_WIRE_807),
	.R_next30(SYNTHESIZED_WIRE_808),
	.R_next31(SYNTHESIZED_WIRE_809),
	.R_next32(SYNTHESIZED_WIRE_810),
	.L_next1(SYNTHESIZED_WIRE_811),
	.L_next2(SYNTHESIZED_WIRE_812),
	.L_next3(SYNTHESIZED_WIRE_813),
	.L_next4(SYNTHESIZED_WIRE_814),
	.L_next5(SYNTHESIZED_WIRE_815),
	.L_next6(SYNTHESIZED_WIRE_816),
	.L_next7(SYNTHESIZED_WIRE_817),
	.L_next8(SYNTHESIZED_WIRE_818),
	.L_next9(SYNTHESIZED_WIRE_819),
	.L_next10(SYNTHESIZED_WIRE_820),
	.L_next11(SYNTHESIZED_WIRE_821),
	.L_next12(SYNTHESIZED_WIRE_822),
	.L_next13(SYNTHESIZED_WIRE_823),
	.L_next14(SYNTHESIZED_WIRE_824),
	.L_next15(SYNTHESIZED_WIRE_825),
	.L_next16(SYNTHESIZED_WIRE_826),
	.L_next17(SYNTHESIZED_WIRE_827),
	.L_next18(SYNTHESIZED_WIRE_828),
	.L_next19(SYNTHESIZED_WIRE_829),
	.L_next20(SYNTHESIZED_WIRE_830),
	.L_next21(SYNTHESIZED_WIRE_831),
	.L_next22(SYNTHESIZED_WIRE_832),
	.L_next23(SYNTHESIZED_WIRE_833),
	.L_next24(SYNTHESIZED_WIRE_834),
	.L_next25(SYNTHESIZED_WIRE_835),
	.L_next26(SYNTHESIZED_WIRE_836),
	.L_next27(SYNTHESIZED_WIRE_837),
	.L_next28(SYNTHESIZED_WIRE_838),
	.L_next29(SYNTHESIZED_WIRE_839),
	.L_next30(SYNTHESIZED_WIRE_840),
	.L_next31(SYNTHESIZED_WIRE_841),
	.L_next32(SYNTHESIZED_WIRE_842));


round	b2v_inst51(
	.R1(SYNTHESIZED_WIRE_779),
	.R2(SYNTHESIZED_WIRE_780),
	.R3(SYNTHESIZED_WIRE_781),
	.R4(SYNTHESIZED_WIRE_782),
	.R5(SYNTHESIZED_WIRE_783),
	.R6(SYNTHESIZED_WIRE_784),
	.R7(SYNTHESIZED_WIRE_785),
	.R8(SYNTHESIZED_WIRE_786),
	.R9(SYNTHESIZED_WIRE_787),
	.R10(SYNTHESIZED_WIRE_788),
	.R11(SYNTHESIZED_WIRE_789),
	.R12(SYNTHESIZED_WIRE_790),
	.R13(SYNTHESIZED_WIRE_791),
	.R14(SYNTHESIZED_WIRE_792),
	.R15(SYNTHESIZED_WIRE_793),
	.R16(SYNTHESIZED_WIRE_794),
	.R17(SYNTHESIZED_WIRE_795),
	.R18(SYNTHESIZED_WIRE_796),
	.R19(SYNTHESIZED_WIRE_797),
	.R20(SYNTHESIZED_WIRE_798),
	.R21(SYNTHESIZED_WIRE_799),
	.R22(SYNTHESIZED_WIRE_800),
	.R23(SYNTHESIZED_WIRE_801),
	.R24(SYNTHESIZED_WIRE_802),
	.R25(SYNTHESIZED_WIRE_803),
	.R26(SYNTHESIZED_WIRE_804),
	.R27(SYNTHESIZED_WIRE_805),
	.R28(SYNTHESIZED_WIRE_806),
	.R29(SYNTHESIZED_WIRE_807),
	.R30(SYNTHESIZED_WIRE_808),
	.R31(SYNTHESIZED_WIRE_809),
	.R32(SYNTHESIZED_WIRE_810),
	.L1(SYNTHESIZED_WIRE_811),
	.L2(SYNTHESIZED_WIRE_812),
	.L3(SYNTHESIZED_WIRE_813),
	.L4(SYNTHESIZED_WIRE_814),
	.L5(SYNTHESIZED_WIRE_815),
	.L6(SYNTHESIZED_WIRE_816),
	.L7(SYNTHESIZED_WIRE_817),
	.L8(SYNTHESIZED_WIRE_818),
	.L9(SYNTHESIZED_WIRE_819),
	.L10(SYNTHESIZED_WIRE_820),
	.L11(SYNTHESIZED_WIRE_821),
	.L12(SYNTHESIZED_WIRE_822),
	.L13(SYNTHESIZED_WIRE_823),
	.L14(SYNTHESIZED_WIRE_824),
	.L15(SYNTHESIZED_WIRE_825),
	.L16(SYNTHESIZED_WIRE_826),
	.L17(SYNTHESIZED_WIRE_827),
	.L18(SYNTHESIZED_WIRE_828),
	.L19(SYNTHESIZED_WIRE_829),
	.L20(SYNTHESIZED_WIRE_830),
	.L21(SYNTHESIZED_WIRE_831),
	.L22(SYNTHESIZED_WIRE_832),
	.L23(SYNTHESIZED_WIRE_833),
	.L24(SYNTHESIZED_WIRE_834),
	.L25(SYNTHESIZED_WIRE_835),
	.L26(SYNTHESIZED_WIRE_836),
	.L27(SYNTHESIZED_WIRE_837),
	.L28(SYNTHESIZED_WIRE_838),
	.L29(SYNTHESIZED_WIRE_839),
	.L30(SYNTHESIZED_WIRE_840),
	.L31(SYNTHESIZED_WIRE_841),
	.L32(SYNTHESIZED_WIRE_842),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_843),
	.R_next1(SYNTHESIZED_WIRE_844),
	.R_next2(SYNTHESIZED_WIRE_845),
	.R_next3(SYNTHESIZED_WIRE_846),
	.R_next4(SYNTHESIZED_WIRE_847),
	.R_next5(SYNTHESIZED_WIRE_848),
	.R_next6(SYNTHESIZED_WIRE_849),
	.R_next7(SYNTHESIZED_WIRE_850),
	.R_next8(SYNTHESIZED_WIRE_851),
	.R_next9(SYNTHESIZED_WIRE_852),
	.R_next10(SYNTHESIZED_WIRE_853),
	.R_next11(SYNTHESIZED_WIRE_854),
	.R_next12(SYNTHESIZED_WIRE_855),
	.R_next13(SYNTHESIZED_WIRE_856),
	.R_next14(SYNTHESIZED_WIRE_857),
	.R_next15(SYNTHESIZED_WIRE_858),
	.R_next16(SYNTHESIZED_WIRE_859),
	.R_next17(SYNTHESIZED_WIRE_860),
	.R_next18(SYNTHESIZED_WIRE_861),
	.R_next19(SYNTHESIZED_WIRE_862),
	.R_next20(SYNTHESIZED_WIRE_863),
	.R_next21(SYNTHESIZED_WIRE_864),
	.R_next22(SYNTHESIZED_WIRE_865),
	.R_next23(SYNTHESIZED_WIRE_866),
	.R_next24(SYNTHESIZED_WIRE_867),
	.R_next25(SYNTHESIZED_WIRE_868),
	.R_next26(SYNTHESIZED_WIRE_869),
	.R_next27(SYNTHESIZED_WIRE_870),
	.R_next28(SYNTHESIZED_WIRE_871),
	.R_next29(SYNTHESIZED_WIRE_872),
	.R_next30(SYNTHESIZED_WIRE_873),
	.R_next31(SYNTHESIZED_WIRE_874),
	.R_next32(SYNTHESIZED_WIRE_875),
	.L_next1(SYNTHESIZED_WIRE_876),
	.L_next2(SYNTHESIZED_WIRE_877),
	.L_next3(SYNTHESIZED_WIRE_878),
	.L_next4(SYNTHESIZED_WIRE_879),
	.L_next5(SYNTHESIZED_WIRE_880),
	.L_next6(SYNTHESIZED_WIRE_881),
	.L_next7(SYNTHESIZED_WIRE_882),
	.L_next8(SYNTHESIZED_WIRE_883),
	.L_next9(SYNTHESIZED_WIRE_884),
	.L_next10(SYNTHESIZED_WIRE_885),
	.L_next11(SYNTHESIZED_WIRE_886),
	.L_next12(SYNTHESIZED_WIRE_887),
	.L_next13(SYNTHESIZED_WIRE_888),
	.L_next14(SYNTHESIZED_WIRE_889),
	.L_next15(SYNTHESIZED_WIRE_890),
	.L_next16(SYNTHESIZED_WIRE_891),
	.L_next17(SYNTHESIZED_WIRE_892),
	.L_next18(SYNTHESIZED_WIRE_893),
	.L_next19(SYNTHESIZED_WIRE_894),
	.L_next20(SYNTHESIZED_WIRE_895),
	.L_next21(SYNTHESIZED_WIRE_896),
	.L_next22(SYNTHESIZED_WIRE_897),
	.L_next23(SYNTHESIZED_WIRE_898),
	.L_next24(SYNTHESIZED_WIRE_899),
	.L_next25(SYNTHESIZED_WIRE_900),
	.L_next26(SYNTHESIZED_WIRE_901),
	.L_next27(SYNTHESIZED_WIRE_902),
	.L_next28(SYNTHESIZED_WIRE_903),
	.L_next29(SYNTHESIZED_WIRE_904),
	.L_next30(SYNTHESIZED_WIRE_905),
	.L_next31(SYNTHESIZED_WIRE_906),
	.L_next32(SYNTHESIZED_WIRE_907));


round	b2v_inst52(
	.R1(SYNTHESIZED_WIRE_844),
	.R2(SYNTHESIZED_WIRE_845),
	.R3(SYNTHESIZED_WIRE_846),
	.R4(SYNTHESIZED_WIRE_847),
	.R5(SYNTHESIZED_WIRE_848),
	.R6(SYNTHESIZED_WIRE_849),
	.R7(SYNTHESIZED_WIRE_850),
	.R8(SYNTHESIZED_WIRE_851),
	.R9(SYNTHESIZED_WIRE_852),
	.R10(SYNTHESIZED_WIRE_853),
	.R11(SYNTHESIZED_WIRE_854),
	.R12(SYNTHESIZED_WIRE_855),
	.R13(SYNTHESIZED_WIRE_856),
	.R14(SYNTHESIZED_WIRE_857),
	.R15(SYNTHESIZED_WIRE_858),
	.R16(SYNTHESIZED_WIRE_859),
	.R17(SYNTHESIZED_WIRE_860),
	.R18(SYNTHESIZED_WIRE_861),
	.R19(SYNTHESIZED_WIRE_862),
	.R20(SYNTHESIZED_WIRE_863),
	.R21(SYNTHESIZED_WIRE_864),
	.R22(SYNTHESIZED_WIRE_865),
	.R23(SYNTHESIZED_WIRE_866),
	.R24(SYNTHESIZED_WIRE_867),
	.R25(SYNTHESIZED_WIRE_868),
	.R26(SYNTHESIZED_WIRE_869),
	.R27(SYNTHESIZED_WIRE_870),
	.R28(SYNTHESIZED_WIRE_871),
	.R29(SYNTHESIZED_WIRE_872),
	.R30(SYNTHESIZED_WIRE_873),
	.R31(SYNTHESIZED_WIRE_874),
	.R32(SYNTHESIZED_WIRE_875),
	.L1(SYNTHESIZED_WIRE_876),
	.L2(SYNTHESIZED_WIRE_877),
	.L3(SYNTHESIZED_WIRE_878),
	.L4(SYNTHESIZED_WIRE_879),
	.L5(SYNTHESIZED_WIRE_880),
	.L6(SYNTHESIZED_WIRE_881),
	.L7(SYNTHESIZED_WIRE_882),
	.L8(SYNTHESIZED_WIRE_883),
	.L9(SYNTHESIZED_WIRE_884),
	.L10(SYNTHESIZED_WIRE_885),
	.L11(SYNTHESIZED_WIRE_886),
	.L12(SYNTHESIZED_WIRE_887),
	.L13(SYNTHESIZED_WIRE_888),
	.L14(SYNTHESIZED_WIRE_889),
	.L15(SYNTHESIZED_WIRE_890),
	.L16(SYNTHESIZED_WIRE_891),
	.L17(SYNTHESIZED_WIRE_892),
	.L18(SYNTHESIZED_WIRE_893),
	.L19(SYNTHESIZED_WIRE_894),
	.L20(SYNTHESIZED_WIRE_895),
	.L21(SYNTHESIZED_WIRE_896),
	.L22(SYNTHESIZED_WIRE_897),
	.L23(SYNTHESIZED_WIRE_898),
	.L24(SYNTHESIZED_WIRE_899),
	.L25(SYNTHESIZED_WIRE_900),
	.L26(SYNTHESIZED_WIRE_901),
	.L27(SYNTHESIZED_WIRE_902),
	.L28(SYNTHESIZED_WIRE_903),
	.L29(SYNTHESIZED_WIRE_904),
	.L30(SYNTHESIZED_WIRE_905),
	.L31(SYNTHESIZED_WIRE_906),
	.L32(SYNTHESIZED_WIRE_907),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_908),
	.R_next1(SYNTHESIZED_WIRE_909),
	.R_next2(SYNTHESIZED_WIRE_910),
	.R_next3(SYNTHESIZED_WIRE_911),
	.R_next4(SYNTHESIZED_WIRE_912),
	.R_next5(SYNTHESIZED_WIRE_913),
	.R_next6(SYNTHESIZED_WIRE_914),
	.R_next7(SYNTHESIZED_WIRE_915),
	.R_next8(SYNTHESIZED_WIRE_916),
	.R_next9(SYNTHESIZED_WIRE_917),
	.R_next10(SYNTHESIZED_WIRE_918),
	.R_next11(SYNTHESIZED_WIRE_919),
	.R_next12(SYNTHESIZED_WIRE_920),
	.R_next13(SYNTHESIZED_WIRE_921),
	.R_next14(SYNTHESIZED_WIRE_922),
	.R_next15(SYNTHESIZED_WIRE_923),
	.R_next16(SYNTHESIZED_WIRE_924),
	.R_next17(SYNTHESIZED_WIRE_925),
	.R_next18(SYNTHESIZED_WIRE_926),
	.R_next19(SYNTHESIZED_WIRE_927),
	.R_next20(SYNTHESIZED_WIRE_928),
	.R_next21(SYNTHESIZED_WIRE_929),
	.R_next22(SYNTHESIZED_WIRE_930),
	.R_next23(SYNTHESIZED_WIRE_931),
	.R_next24(SYNTHESIZED_WIRE_932),
	.R_next25(SYNTHESIZED_WIRE_933),
	.R_next26(SYNTHESIZED_WIRE_934),
	.R_next27(SYNTHESIZED_WIRE_935),
	.R_next28(SYNTHESIZED_WIRE_936),
	.R_next29(SYNTHESIZED_WIRE_937),
	.R_next30(SYNTHESIZED_WIRE_938),
	.R_next31(SYNTHESIZED_WIRE_939),
	.R_next32(SYNTHESIZED_WIRE_940),
	.L_next1(SYNTHESIZED_WIRE_941),
	.L_next2(SYNTHESIZED_WIRE_942),
	.L_next3(SYNTHESIZED_WIRE_943),
	.L_next4(SYNTHESIZED_WIRE_944),
	.L_next5(SYNTHESIZED_WIRE_945),
	.L_next6(SYNTHESIZED_WIRE_946),
	.L_next7(SYNTHESIZED_WIRE_947),
	.L_next8(SYNTHESIZED_WIRE_948),
	.L_next9(SYNTHESIZED_WIRE_949),
	.L_next10(SYNTHESIZED_WIRE_950),
	.L_next11(SYNTHESIZED_WIRE_951),
	.L_next12(SYNTHESIZED_WIRE_952),
	.L_next13(SYNTHESIZED_WIRE_953),
	.L_next14(SYNTHESIZED_WIRE_954),
	.L_next15(SYNTHESIZED_WIRE_955),
	.L_next16(SYNTHESIZED_WIRE_956),
	.L_next17(SYNTHESIZED_WIRE_957),
	.L_next18(SYNTHESIZED_WIRE_958),
	.L_next19(SYNTHESIZED_WIRE_959),
	.L_next20(SYNTHESIZED_WIRE_960),
	.L_next21(SYNTHESIZED_WIRE_961),
	.L_next22(SYNTHESIZED_WIRE_962),
	.L_next23(SYNTHESIZED_WIRE_963),
	.L_next24(SYNTHESIZED_WIRE_964),
	.L_next25(SYNTHESIZED_WIRE_965),
	.L_next26(SYNTHESIZED_WIRE_966),
	.L_next27(SYNTHESIZED_WIRE_967),
	.L_next28(SYNTHESIZED_WIRE_968),
	.L_next29(SYNTHESIZED_WIRE_969),
	.L_next30(SYNTHESIZED_WIRE_970),
	.L_next31(SYNTHESIZED_WIRE_971),
	.L_next32(SYNTHESIZED_WIRE_972));


round	b2v_inst53(
	.R1(SYNTHESIZED_WIRE_909),
	.R2(SYNTHESIZED_WIRE_910),
	.R3(SYNTHESIZED_WIRE_911),
	.R4(SYNTHESIZED_WIRE_912),
	.R5(SYNTHESIZED_WIRE_913),
	.R6(SYNTHESIZED_WIRE_914),
	.R7(SYNTHESIZED_WIRE_915),
	.R8(SYNTHESIZED_WIRE_916),
	.R9(SYNTHESIZED_WIRE_917),
	.R10(SYNTHESIZED_WIRE_918),
	.R11(SYNTHESIZED_WIRE_919),
	.R12(SYNTHESIZED_WIRE_920),
	.R13(SYNTHESIZED_WIRE_921),
	.R14(SYNTHESIZED_WIRE_922),
	.R15(SYNTHESIZED_WIRE_923),
	.R16(SYNTHESIZED_WIRE_924),
	.R17(SYNTHESIZED_WIRE_925),
	.R18(SYNTHESIZED_WIRE_926),
	.R19(SYNTHESIZED_WIRE_927),
	.R20(SYNTHESIZED_WIRE_928),
	.R21(SYNTHESIZED_WIRE_929),
	.R22(SYNTHESIZED_WIRE_930),
	.R23(SYNTHESIZED_WIRE_931),
	.R24(SYNTHESIZED_WIRE_932),
	.R25(SYNTHESIZED_WIRE_933),
	.R26(SYNTHESIZED_WIRE_934),
	.R27(SYNTHESIZED_WIRE_935),
	.R28(SYNTHESIZED_WIRE_936),
	.R29(SYNTHESIZED_WIRE_937),
	.R30(SYNTHESIZED_WIRE_938),
	.R31(SYNTHESIZED_WIRE_939),
	.R32(SYNTHESIZED_WIRE_940),
	.L1(SYNTHESIZED_WIRE_941),
	.L2(SYNTHESIZED_WIRE_942),
	.L3(SYNTHESIZED_WIRE_943),
	.L4(SYNTHESIZED_WIRE_944),
	.L5(SYNTHESIZED_WIRE_945),
	.L6(SYNTHESIZED_WIRE_946),
	.L7(SYNTHESIZED_WIRE_947),
	.L8(SYNTHESIZED_WIRE_948),
	.L9(SYNTHESIZED_WIRE_949),
	.L10(SYNTHESIZED_WIRE_950),
	.L11(SYNTHESIZED_WIRE_951),
	.L12(SYNTHESIZED_WIRE_952),
	.L13(SYNTHESIZED_WIRE_953),
	.L14(SYNTHESIZED_WIRE_954),
	.L15(SYNTHESIZED_WIRE_955),
	.L16(SYNTHESIZED_WIRE_956),
	.L17(SYNTHESIZED_WIRE_957),
	.L18(SYNTHESIZED_WIRE_958),
	.L19(SYNTHESIZED_WIRE_959),
	.L20(SYNTHESIZED_WIRE_960),
	.L21(SYNTHESIZED_WIRE_961),
	.L22(SYNTHESIZED_WIRE_962),
	.L23(SYNTHESIZED_WIRE_963),
	.L24(SYNTHESIZED_WIRE_964),
	.L25(SYNTHESIZED_WIRE_965),
	.L26(SYNTHESIZED_WIRE_966),
	.L27(SYNTHESIZED_WIRE_967),
	.L28(SYNTHESIZED_WIRE_968),
	.L29(SYNTHESIZED_WIRE_969),
	.L30(SYNTHESIZED_WIRE_970),
	.L31(SYNTHESIZED_WIRE_971),
	.L32(SYNTHESIZED_WIRE_972),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_973),
	.R_next1(SYNTHESIZED_WIRE_974),
	.R_next2(SYNTHESIZED_WIRE_975),
	.R_next3(SYNTHESIZED_WIRE_976),
	.R_next4(SYNTHESIZED_WIRE_977),
	.R_next5(SYNTHESIZED_WIRE_978),
	.R_next6(SYNTHESIZED_WIRE_979),
	.R_next7(SYNTHESIZED_WIRE_980),
	.R_next8(SYNTHESIZED_WIRE_981),
	.R_next9(SYNTHESIZED_WIRE_982),
	.R_next10(SYNTHESIZED_WIRE_983),
	.R_next11(SYNTHESIZED_WIRE_984),
	.R_next12(SYNTHESIZED_WIRE_985),
	.R_next13(SYNTHESIZED_WIRE_986),
	.R_next14(SYNTHESIZED_WIRE_987),
	.R_next15(SYNTHESIZED_WIRE_988),
	.R_next16(SYNTHESIZED_WIRE_989),
	.R_next17(SYNTHESIZED_WIRE_990),
	.R_next18(SYNTHESIZED_WIRE_991),
	.R_next19(SYNTHESIZED_WIRE_992),
	.R_next20(SYNTHESIZED_WIRE_993),
	.R_next21(SYNTHESIZED_WIRE_994),
	.R_next22(SYNTHESIZED_WIRE_995),
	.R_next23(SYNTHESIZED_WIRE_996),
	.R_next24(SYNTHESIZED_WIRE_997),
	.R_next25(SYNTHESIZED_WIRE_998),
	.R_next26(SYNTHESIZED_WIRE_999),
	.R_next27(SYNTHESIZED_WIRE_1000),
	.R_next28(SYNTHESIZED_WIRE_1001),
	.R_next29(SYNTHESIZED_WIRE_1002),
	.R_next30(SYNTHESIZED_WIRE_1003),
	.R_next31(SYNTHESIZED_WIRE_1004),
	.R_next32(SYNTHESIZED_WIRE_1005),
	.L_next1(SYNTHESIZED_WIRE_1006),
	.L_next2(SYNTHESIZED_WIRE_1007),
	.L_next3(SYNTHESIZED_WIRE_1008),
	.L_next4(SYNTHESIZED_WIRE_1009),
	.L_next5(SYNTHESIZED_WIRE_1010),
	.L_next6(SYNTHESIZED_WIRE_1011),
	.L_next7(SYNTHESIZED_WIRE_1012),
	.L_next8(SYNTHESIZED_WIRE_1013),
	.L_next9(SYNTHESIZED_WIRE_1014),
	.L_next10(SYNTHESIZED_WIRE_1015),
	.L_next11(SYNTHESIZED_WIRE_1016),
	.L_next12(SYNTHESIZED_WIRE_1017),
	.L_next13(SYNTHESIZED_WIRE_1018),
	.L_next14(SYNTHESIZED_WIRE_1019),
	.L_next15(SYNTHESIZED_WIRE_1020),
	.L_next16(SYNTHESIZED_WIRE_1021),
	.L_next17(SYNTHESIZED_WIRE_1022),
	.L_next18(SYNTHESIZED_WIRE_1023),
	.L_next19(SYNTHESIZED_WIRE_1024),
	.L_next20(SYNTHESIZED_WIRE_1025),
	.L_next21(SYNTHESIZED_WIRE_1026),
	.L_next22(SYNTHESIZED_WIRE_1027),
	.L_next23(SYNTHESIZED_WIRE_1028),
	.L_next24(SYNTHESIZED_WIRE_1029),
	.L_next25(SYNTHESIZED_WIRE_1030),
	.L_next26(SYNTHESIZED_WIRE_1031),
	.L_next27(SYNTHESIZED_WIRE_1032),
	.L_next28(SYNTHESIZED_WIRE_1033),
	.L_next29(SYNTHESIZED_WIRE_1034),
	.L_next30(SYNTHESIZED_WIRE_1035),
	.L_next31(SYNTHESIZED_WIRE_1036),
	.L_next32(SYNTHESIZED_WIRE_1037));


round	b2v_inst54(
	.R1(SYNTHESIZED_WIRE_974),
	.R2(SYNTHESIZED_WIRE_975),
	.R3(SYNTHESIZED_WIRE_976),
	.R4(SYNTHESIZED_WIRE_977),
	.R5(SYNTHESIZED_WIRE_978),
	.R6(SYNTHESIZED_WIRE_979),
	.R7(SYNTHESIZED_WIRE_980),
	.R8(SYNTHESIZED_WIRE_981),
	.R9(SYNTHESIZED_WIRE_982),
	.R10(SYNTHESIZED_WIRE_983),
	.R11(SYNTHESIZED_WIRE_984),
	.R12(SYNTHESIZED_WIRE_985),
	.R13(SYNTHESIZED_WIRE_986),
	.R14(SYNTHESIZED_WIRE_987),
	.R15(SYNTHESIZED_WIRE_988),
	.R16(SYNTHESIZED_WIRE_989),
	.R17(SYNTHESIZED_WIRE_990),
	.R18(SYNTHESIZED_WIRE_991),
	.R19(SYNTHESIZED_WIRE_992),
	.R20(SYNTHESIZED_WIRE_993),
	.R21(SYNTHESIZED_WIRE_994),
	.R22(SYNTHESIZED_WIRE_995),
	.R23(SYNTHESIZED_WIRE_996),
	.R24(SYNTHESIZED_WIRE_997),
	.R25(SYNTHESIZED_WIRE_998),
	.R26(SYNTHESIZED_WIRE_999),
	.R27(SYNTHESIZED_WIRE_1000),
	.R28(SYNTHESIZED_WIRE_1001),
	.R29(SYNTHESIZED_WIRE_1002),
	.R30(SYNTHESIZED_WIRE_1003),
	.R31(SYNTHESIZED_WIRE_1004),
	.R32(SYNTHESIZED_WIRE_1005),
	.L1(SYNTHESIZED_WIRE_1006),
	.L2(SYNTHESIZED_WIRE_1007),
	.L3(SYNTHESIZED_WIRE_1008),
	.L4(SYNTHESIZED_WIRE_1009),
	.L5(SYNTHESIZED_WIRE_1010),
	.L6(SYNTHESIZED_WIRE_1011),
	.L7(SYNTHESIZED_WIRE_1012),
	.L8(SYNTHESIZED_WIRE_1013),
	.L9(SYNTHESIZED_WIRE_1014),
	.L10(SYNTHESIZED_WIRE_1015),
	.L11(SYNTHESIZED_WIRE_1016),
	.L12(SYNTHESIZED_WIRE_1017),
	.L13(SYNTHESIZED_WIRE_1018),
	.L14(SYNTHESIZED_WIRE_1019),
	.L15(SYNTHESIZED_WIRE_1020),
	.L16(SYNTHESIZED_WIRE_1021),
	.L17(SYNTHESIZED_WIRE_1022),
	.L18(SYNTHESIZED_WIRE_1023),
	.L19(SYNTHESIZED_WIRE_1024),
	.L20(SYNTHESIZED_WIRE_1025),
	.L21(SYNTHESIZED_WIRE_1026),
	.L22(SYNTHESIZED_WIRE_1027),
	.L23(SYNTHESIZED_WIRE_1028),
	.L24(SYNTHESIZED_WIRE_1029),
	.L25(SYNTHESIZED_WIRE_1030),
	.L26(SYNTHESIZED_WIRE_1031),
	.L27(SYNTHESIZED_WIRE_1032),
	.L28(SYNTHESIZED_WIRE_1033),
	.L29(SYNTHESIZED_WIRE_1034),
	.L30(SYNTHESIZED_WIRE_1035),
	.L31(SYNTHESIZED_WIRE_1036),
	.L32(SYNTHESIZED_WIRE_1037),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_1038),
	.R_next1(SYNTHESIZED_WIRE_1039),
	.R_next2(SYNTHESIZED_WIRE_1040),
	.R_next3(SYNTHESIZED_WIRE_1041),
	.R_next4(SYNTHESIZED_WIRE_1042),
	.R_next5(SYNTHESIZED_WIRE_1043),
	.R_next6(SYNTHESIZED_WIRE_1044),
	.R_next7(SYNTHESIZED_WIRE_1045),
	.R_next8(SYNTHESIZED_WIRE_1046),
	.R_next9(SYNTHESIZED_WIRE_1047),
	.R_next10(SYNTHESIZED_WIRE_1048),
	.R_next11(SYNTHESIZED_WIRE_1049),
	.R_next12(SYNTHESIZED_WIRE_1050),
	.R_next13(SYNTHESIZED_WIRE_1051),
	.R_next14(SYNTHESIZED_WIRE_1052),
	.R_next15(SYNTHESIZED_WIRE_1053),
	.R_next16(SYNTHESIZED_WIRE_1054),
	.R_next17(SYNTHESIZED_WIRE_1055),
	.R_next18(SYNTHESIZED_WIRE_1056),
	.R_next19(SYNTHESIZED_WIRE_1057),
	.R_next20(SYNTHESIZED_WIRE_1058),
	.R_next21(SYNTHESIZED_WIRE_1059),
	.R_next22(SYNTHESIZED_WIRE_1060),
	.R_next23(SYNTHESIZED_WIRE_1061),
	.R_next24(SYNTHESIZED_WIRE_1062),
	.R_next25(SYNTHESIZED_WIRE_1063),
	.R_next26(SYNTHESIZED_WIRE_1064),
	.R_next27(SYNTHESIZED_WIRE_1065),
	.R_next28(SYNTHESIZED_WIRE_1066),
	.R_next29(SYNTHESIZED_WIRE_1067),
	.R_next30(SYNTHESIZED_WIRE_1068),
	.R_next31(SYNTHESIZED_WIRE_1069),
	.R_next32(SYNTHESIZED_WIRE_1070),
	.L_next1(SYNTHESIZED_WIRE_1071),
	.L_next2(SYNTHESIZED_WIRE_1072),
	.L_next3(SYNTHESIZED_WIRE_1073),
	.L_next4(SYNTHESIZED_WIRE_1074),
	.L_next5(SYNTHESIZED_WIRE_1075),
	.L_next6(SYNTHESIZED_WIRE_1076),
	.L_next7(SYNTHESIZED_WIRE_1077),
	.L_next8(SYNTHESIZED_WIRE_1078),
	.L_next9(SYNTHESIZED_WIRE_1079),
	.L_next10(SYNTHESIZED_WIRE_1080),
	.L_next11(SYNTHESIZED_WIRE_1081),
	.L_next12(SYNTHESIZED_WIRE_1082),
	.L_next13(SYNTHESIZED_WIRE_1083),
	.L_next14(SYNTHESIZED_WIRE_1084),
	.L_next15(SYNTHESIZED_WIRE_1085),
	.L_next16(SYNTHESIZED_WIRE_1086),
	.L_next17(SYNTHESIZED_WIRE_1087),
	.L_next18(SYNTHESIZED_WIRE_1088),
	.L_next19(SYNTHESIZED_WIRE_1089),
	.L_next20(SYNTHESIZED_WIRE_1090),
	.L_next21(SYNTHESIZED_WIRE_1091),
	.L_next22(SYNTHESIZED_WIRE_1092),
	.L_next23(SYNTHESIZED_WIRE_1093),
	.L_next24(SYNTHESIZED_WIRE_1094),
	.L_next25(SYNTHESIZED_WIRE_1095),
	.L_next26(SYNTHESIZED_WIRE_1096),
	.L_next27(SYNTHESIZED_WIRE_1097),
	.L_next28(SYNTHESIZED_WIRE_1098),
	.L_next29(SYNTHESIZED_WIRE_1099),
	.L_next30(SYNTHESIZED_WIRE_1100),
	.L_next31(SYNTHESIZED_WIRE_1101),
	.L_next32(SYNTHESIZED_WIRE_1102));


round	b2v_inst55(
	.R1(SYNTHESIZED_WIRE_1039),
	.R2(SYNTHESIZED_WIRE_1040),
	.R3(SYNTHESIZED_WIRE_1041),
	.R4(SYNTHESIZED_WIRE_1042),
	.R5(SYNTHESIZED_WIRE_1043),
	.R6(SYNTHESIZED_WIRE_1044),
	.R7(SYNTHESIZED_WIRE_1045),
	.R8(SYNTHESIZED_WIRE_1046),
	.R9(SYNTHESIZED_WIRE_1047),
	.R10(SYNTHESIZED_WIRE_1048),
	.R11(SYNTHESIZED_WIRE_1049),
	.R12(SYNTHESIZED_WIRE_1050),
	.R13(SYNTHESIZED_WIRE_1051),
	.R14(SYNTHESIZED_WIRE_1052),
	.R15(SYNTHESIZED_WIRE_1053),
	.R16(SYNTHESIZED_WIRE_1054),
	.R17(SYNTHESIZED_WIRE_1055),
	.R18(SYNTHESIZED_WIRE_1056),
	.R19(SYNTHESIZED_WIRE_1057),
	.R20(SYNTHESIZED_WIRE_1058),
	.R21(SYNTHESIZED_WIRE_1059),
	.R22(SYNTHESIZED_WIRE_1060),
	.R23(SYNTHESIZED_WIRE_1061),
	.R24(SYNTHESIZED_WIRE_1062),
	.R25(SYNTHESIZED_WIRE_1063),
	.R26(SYNTHESIZED_WIRE_1064),
	.R27(SYNTHESIZED_WIRE_1065),
	.R28(SYNTHESIZED_WIRE_1066),
	.R29(SYNTHESIZED_WIRE_1067),
	.R30(SYNTHESIZED_WIRE_1068),
	.R31(SYNTHESIZED_WIRE_1069),
	.R32(SYNTHESIZED_WIRE_1070),
	.L1(SYNTHESIZED_WIRE_1071),
	.L2(SYNTHESIZED_WIRE_1072),
	.L3(SYNTHESIZED_WIRE_1073),
	.L4(SYNTHESIZED_WIRE_1074),
	.L5(SYNTHESIZED_WIRE_1075),
	.L6(SYNTHESIZED_WIRE_1076),
	.L7(SYNTHESIZED_WIRE_1077),
	.L8(SYNTHESIZED_WIRE_1078),
	.L9(SYNTHESIZED_WIRE_1079),
	.L10(SYNTHESIZED_WIRE_1080),
	.L11(SYNTHESIZED_WIRE_1081),
	.L12(SYNTHESIZED_WIRE_1082),
	.L13(SYNTHESIZED_WIRE_1083),
	.L14(SYNTHESIZED_WIRE_1084),
	.L15(SYNTHESIZED_WIRE_1085),
	.L16(SYNTHESIZED_WIRE_1086),
	.L17(SYNTHESIZED_WIRE_1087),
	.L18(SYNTHESIZED_WIRE_1088),
	.L19(SYNTHESIZED_WIRE_1089),
	.L20(SYNTHESIZED_WIRE_1090),
	.L21(SYNTHESIZED_WIRE_1091),
	.L22(SYNTHESIZED_WIRE_1092),
	.L23(SYNTHESIZED_WIRE_1093),
	.L24(SYNTHESIZED_WIRE_1094),
	.L25(SYNTHESIZED_WIRE_1095),
	.L26(SYNTHESIZED_WIRE_1096),
	.L27(SYNTHESIZED_WIRE_1097),
	.L28(SYNTHESIZED_WIRE_1098),
	.L29(SYNTHESIZED_WIRE_1099),
	.L30(SYNTHESIZED_WIRE_1100),
	.L31(SYNTHESIZED_WIRE_1101),
	.L32(SYNTHESIZED_WIRE_1102),
	.clk(clk),
	.rst_n(rst_n),
	.key(SYNTHESIZED_WIRE_1103),
	.R_next1(SYNTHESIZED_WIRE_195),
	.R_next2(SYNTHESIZED_WIRE_196),
	.R_next3(SYNTHESIZED_WIRE_197),
	.R_next4(SYNTHESIZED_WIRE_198),
	.R_next5(SYNTHESIZED_WIRE_199),
	.R_next6(SYNTHESIZED_WIRE_200),
	.R_next7(SYNTHESIZED_WIRE_201),
	.R_next8(SYNTHESIZED_WIRE_202),
	.R_next9(SYNTHESIZED_WIRE_203),
	.R_next10(SYNTHESIZED_WIRE_204),
	.R_next11(SYNTHESIZED_WIRE_205),
	.R_next12(SYNTHESIZED_WIRE_206),
	.R_next13(SYNTHESIZED_WIRE_207),
	.R_next14(SYNTHESIZED_WIRE_208),
	.R_next15(SYNTHESIZED_WIRE_209),
	.R_next16(SYNTHESIZED_WIRE_210),
	.R_next17(SYNTHESIZED_WIRE_211),
	.R_next18(SYNTHESIZED_WIRE_212),
	.R_next19(SYNTHESIZED_WIRE_213),
	.R_next20(SYNTHESIZED_WIRE_214),
	.R_next21(SYNTHESIZED_WIRE_215),
	.R_next22(SYNTHESIZED_WIRE_216),
	.R_next23(SYNTHESIZED_WIRE_217),
	.R_next24(SYNTHESIZED_WIRE_218),
	.R_next25(SYNTHESIZED_WIRE_219),
	.R_next26(SYNTHESIZED_WIRE_220),
	.R_next27(SYNTHESIZED_WIRE_221),
	.R_next28(SYNTHESIZED_WIRE_222),
	.R_next29(SYNTHESIZED_WIRE_223),
	.R_next30(SYNTHESIZED_WIRE_224),
	.R_next31(SYNTHESIZED_WIRE_225),
	.R_next32(SYNTHESIZED_WIRE_226),
	.L_next1(SYNTHESIZED_WIRE_227),
	.L_next2(SYNTHESIZED_WIRE_228),
	.L_next3(SYNTHESIZED_WIRE_229),
	.L_next4(SYNTHESIZED_WIRE_230),
	.L_next5(SYNTHESIZED_WIRE_231),
	.L_next6(SYNTHESIZED_WIRE_232),
	.L_next7(SYNTHESIZED_WIRE_233),
	.L_next8(SYNTHESIZED_WIRE_234),
	.L_next9(SYNTHESIZED_WIRE_235),
	.L_next10(SYNTHESIZED_WIRE_236),
	.L_next11(SYNTHESIZED_WIRE_237),
	.L_next12(SYNTHESIZED_WIRE_238),
	.L_next13(SYNTHESIZED_WIRE_239),
	.L_next14(SYNTHESIZED_WIRE_240),
	.L_next15(SYNTHESIZED_WIRE_241),
	.L_next16(SYNTHESIZED_WIRE_242),
	.L_next17(SYNTHESIZED_WIRE_243),
	.L_next18(SYNTHESIZED_WIRE_244),
	.L_next19(SYNTHESIZED_WIRE_245),
	.L_next20(SYNTHESIZED_WIRE_246),
	.L_next21(SYNTHESIZED_WIRE_247),
	.L_next22(SYNTHESIZED_WIRE_248),
	.L_next23(SYNTHESIZED_WIRE_249),
	.L_next24(SYNTHESIZED_WIRE_250),
	.L_next25(SYNTHESIZED_WIRE_251),
	.L_next26(SYNTHESIZED_WIRE_252),
	.L_next27(SYNTHESIZED_WIRE_253),
	.L_next28(SYNTHESIZED_WIRE_254),
	.L_next29(SYNTHESIZED_WIRE_255),
	.L_next30(SYNTHESIZED_WIRE_256),
	.L_next31(SYNTHESIZED_WIRE_257),
	.L_next32(SYNTHESIZED_WIRE_258));

assign	des_encrypt_out = des_encrypt_out_ALTERA_SYNTHESIZED;

endmodule
