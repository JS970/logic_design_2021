// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Nov 24 22:19:19 2021"

module lshift2(
	in14,
	in28,
	in27,
	in26,
	in25,
	in24,
	in23,
	in22,
	in21,
	in20,
	in19,
	in18,
	in17,
	in16,
	in15,
	in13,
	in12,
	in11,
	in10,
	in9,
	in8,
	in7,
	in6,
	in5,
	in4,
	in3,
	in2,
	in1,
	out28,
	out27,
	out26,
	out25,
	out24,
	out23,
	out22,
	out21,
	out20,
	out19,
	out18,
	out17,
	out16,
	out15,
	out14,
	out13,
	out12,
	out11,
	out10,
	out9,
	out8,
	out7,
	out6,
	out5,
	out4,
	out3,
	out2,
	out1
);


input wire	in14;
input wire	in28;
input wire	in27;
input wire	in26;
input wire	in25;
input wire	in24;
input wire	in23;
input wire	in22;
input wire	in21;
input wire	in20;
input wire	in19;
input wire	in18;
input wire	in17;
input wire	in16;
input wire	in15;
input wire	in13;
input wire	in12;
input wire	in11;
input wire	in10;
input wire	in9;
input wire	in8;
input wire	in7;
input wire	in6;
input wire	in5;
input wire	in4;
input wire	in3;
input wire	in2;
input wire	in1;
output wire	out28;
output wire	out27;
output wire	out26;
output wire	out25;
output wire	out24;
output wire	out23;
output wire	out22;
output wire	out21;
output wire	out20;
output wire	out19;
output wire	out18;
output wire	out17;
output wire	out16;
output wire	out15;
output wire	out14;
output wire	out13;
output wire	out12;
output wire	out11;
output wire	out10;
output wire	out9;
output wire	out8;
output wire	out7;
output wire	out6;
output wire	out5;
output wire	out4;
output wire	out3;
output wire	out2;
output wire	out1;


assign	out28 = in26;
assign	out27 = in25;
assign	out26 = in24;
assign	out25 = in23;
assign	out24 = in22;
assign	out23 = in21;
assign	out22 = in20;
assign	out21 = in19;
assign	out20 = in18;
assign	out19 = in17;
assign	out18 = in16;
assign	out17 = in15;
assign	out16 = in14;
assign	out15 = in13;
assign	out14 = in12;
assign	out13 = in11;
assign	out12 = in10;
assign	out11 = in9;
assign	out10 = in8;
assign	out9 = in7;
assign	out8 = in6;
assign	out7 = in5;
assign	out6 = in4;
assign	out5 = in3;
assign	out4 = in2;
assign	out3 = in1;
assign	out2 = in28;
assign	out1 = in27;




endmodule
