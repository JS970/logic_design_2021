// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Sat Nov 20 17:40:51 2021"

module b2seg_bus(
	b_in,
	a,
	b,
	c,
	d,
	e,
	f,
	g
);


input wire	[3:0] b_in;
output wire	a;
output wire	b;
output wire	c;
output wire	d;
output wire	e;
output wire	f;
output wire	g;

wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_144;

assign	SYNTHESIZED_WIRE_144 = 0;



assign	SYNTHESIZED_WIRE_143 =  ~b_in[3];

assign	SYNTHESIZED_WIRE_124 =  ~b_in[2];

assign	SYNTHESIZED_WIRE_128 = b_in[3] & SYNTHESIZED_WIRE_124 & b_in[1] & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_127 = b_in[3] & b_in[2] & b_in[1] & b_in[0];

assign	SYNTHESIZED_WIRE_129 = b_in[3] & b_in[2] & b_in[1] & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_130 = b_in[3] & b_in[2] & SYNTHESIZED_WIRE_126 & b_in[0];

assign	SYNTHESIZED_WIRE_132 = b_in[3] & b_in[2] & SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_131 = b_in[3] & SYNTHESIZED_WIRE_124 & b_in[1] & b_in[0];

assign	SYNTHESIZED_WIRE_126 =  ~b_in[1];

assign	SYNTHESIZED_WIRE_125 =  ~b_in[0];

assign	a = SYNTHESIZED_WIRE_127 | SYNTHESIZED_WIRE_128 | SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_129;

assign	b = SYNTHESIZED_WIRE_129 | SYNTHESIZED_WIRE_128 | SYNTHESIZED_WIRE_13 | SYNTHESIZED_WIRE_130;

assign	c = SYNTHESIZED_WIRE_131 | SYNTHESIZED_WIRE_128 | SYNTHESIZED_WIRE_17 | SYNTHESIZED_WIRE_130;

assign	f = SYNTHESIZED_WIRE_127 | SYNTHESIZED_WIRE_131 | SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_129;

assign	d = SYNTHESIZED_WIRE_129 | SYNTHESIZED_WIRE_132 | SYNTHESIZED_WIRE_130 | SYNTHESIZED_WIRE_131 | SYNTHESIZED_WIRE_128 | SYNTHESIZED_WIRE_28;

assign	SYNTHESIZED_WIRE_42 = SYNTHESIZED_WIRE_127 | SYNTHESIZED_WIRE_130 | SYNTHESIZED_WIRE_129 | SYNTHESIZED_WIRE_132 | SYNTHESIZED_WIRE_131 | SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_44 = SYNTHESIZED_WIRE_127 | SYNTHESIZED_WIRE_130 | SYNTHESIZED_WIRE_129 | SYNTHESIZED_WIRE_132 | SYNTHESIZED_WIRE_131 | SYNTHESIZED_WIRE_128;

assign	e = SYNTHESIZED_WIRE_41 | SYNTHESIZED_WIRE_42;

assign	g = SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_140 = b_in[3] & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_126 & b_in[0];

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_134 | SYNTHESIZED_WIRE_135 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_137 | SYNTHESIZED_WIRE_138 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_140;

assign	SYNTHESIZED_WIRE_139 = b_in[3] & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_135 | SYNTHESIZED_WIRE_138 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_142 | SYNTHESIZED_WIRE_137 | SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_137 = SYNTHESIZED_WIRE_143 & b_in[2] & b_in[1] & b_in[0];

assign	SYNTHESIZED_WIRE_141 = SYNTHESIZED_WIRE_125 & SYNTHESIZED_WIRE_143 & b_in[2] & b_in[1];

assign	SYNTHESIZED_WIRE_142 = SYNTHESIZED_WIRE_143 & b_in[2] & SYNTHESIZED_WIRE_126 & b_in[0];

assign	SYNTHESIZED_WIRE_28 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_134 | SYNTHESIZED_WIRE_142 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_140 | SYNTHESIZED_WIRE_144;

assign	SYNTHESIZED_WIRE_138 = SYNTHESIZED_WIRE_143 & b_in[2] & SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_136 = SYNTHESIZED_WIRE_143 & SYNTHESIZED_WIRE_124 & b_in[1] & b_in[0];

assign	SYNTHESIZED_WIRE_134 = SYNTHESIZED_WIRE_143 & SYNTHESIZED_WIRE_124 & b_in[1] & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_135 = SYNTHESIZED_WIRE_143 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_126 & b_in[0];

assign	SYNTHESIZED_WIRE_133 = SYNTHESIZED_WIRE_143 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_134 | SYNTHESIZED_WIRE_142 | SYNTHESIZED_WIRE_137 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_140;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_142 | SYNTHESIZED_WIRE_138 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_137 | SYNTHESIZED_WIRE_140 | SYNTHESIZED_WIRE_144;

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_140 | SYNTHESIZED_WIRE_139;

assign	SYNTHESIZED_WIRE_41 = SYNTHESIZED_WIRE_133 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_134;

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_134 | SYNTHESIZED_WIRE_138 | SYNTHESIZED_WIRE_136 | SYNTHESIZED_WIRE_142 | SYNTHESIZED_WIRE_139 | SYNTHESIZED_WIRE_141 | SYNTHESIZED_WIRE_140 | SYNTHESIZED_WIRE_144;



endmodule
