// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Nov 24 20:45:44 2021"

module s_box_6(
	clk,
	rst_n,
	sbox1_in,
	sbox1_out
);


input wire	clk;
input wire	rst_n;
input wire	[5:0] sbox1_in;
output wire	[3:0] sbox1_out;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	[3:0] SYNTHESIZED_WIRE_12;
wire	[3:0] SYNTHESIZED_WIRE_13;
wire	[3:0] SYNTHESIZED_WIRE_14;
wire	[3:0] SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	[3:0] SYNTHESIZED_WIRE_17;
wire	[3:0] SYNTHESIZED_WIRE_18;
wire	[3:0] SYNTHESIZED_WIRE_19;
wire	[3:0] SYNTHESIZED_WIRE_20;
wire	[3:0] SYNTHESIZED_WIRE_21;
wire	[3:0] SYNTHESIZED_WIRE_22;
wire	[3:0] SYNTHESIZED_WIRE_23;
wire	[3:0] SYNTHESIZED_WIRE_24;
wire	[3:0] SYNTHESIZED_WIRE_25;
wire	[3:0] SYNTHESIZED_WIRE_26;
wire	[3:0] SYNTHESIZED_WIRE_27;
wire	[3:0] SYNTHESIZED_WIRE_28;
wire	[3:0] SYNTHESIZED_WIRE_29;
wire	[3:0] SYNTHESIZED_WIRE_30;
wire	[3:0] SYNTHESIZED_WIRE_31;
wire	[3:0] SYNTHESIZED_WIRE_32;
wire	[3:0] SYNTHESIZED_WIRE_33;
wire	[3:0] SYNTHESIZED_WIRE_34;
wire	[3:0] SYNTHESIZED_WIRE_35;
wire	[3:0] SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	[3:0] SYNTHESIZED_WIRE_38;
wire	[3:0] SYNTHESIZED_WIRE_39;
wire	[3:0] SYNTHESIZED_WIRE_40;
wire	[3:0] SYNTHESIZED_WIRE_41;
wire	[3:0] SYNTHESIZED_WIRE_42;
wire	[3:0] SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_71;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;





six_bit_decoder	b2v_inst(
	.Din(sbox1_in),
	.D1(SYNTHESIZED_WIRE_93),
	.D2(SYNTHESIZED_WIRE_85),
	.D3(SYNTHESIZED_WIRE_52),
	.D4(SYNTHESIZED_WIRE_101),
	.D5(SYNTHESIZED_WIRE_88),
	.D6(SYNTHESIZED_WIRE_0),
	.D7(SYNTHESIZED_WIRE_104),
	.D8(SYNTHESIZED_WIRE_56),
	.D9(SYNTHESIZED_WIRE_81),
	.D10(SYNTHESIZED_WIRE_73),
	.D11(SYNTHESIZED_WIRE_59),
	.D12(SYNTHESIZED_WIRE_96),
	.D13(SYNTHESIZED_WIRE_68),
	.D14(SYNTHESIZED_WIRE_84),
	.D15(SYNTHESIZED_WIRE_77),
	.D16(SYNTHESIZED_WIRE_64),
	.D17(SYNTHESIZED_WIRE_48),
	.D18(SYNTHESIZED_WIRE_71),
	.D19(SYNTHESIZED_WIRE_97),
	.D20(SYNTHESIZED_WIRE_55),
	.D21(SYNTHESIZED_WIRE_60),
	.D22(SYNTHESIZED_WIRE_100),
	.D23(SYNTHESIZED_WIRE_3),
	.D24(SYNTHESIZED_WIRE_44),
	.D25(SYNTHESIZED_WIRE_47),
	.D26(SYNTHESIZED_WIRE_51),
	.D27(SYNTHESIZED_WIRE_76),
	.D28(SYNTHESIZED_WIRE_89),
	.D29(SYNTHESIZED_WIRE_67),
	.D30(SYNTHESIZED_WIRE_63),
	.D31(SYNTHESIZED_WIRE_92),
	.D32(SYNTHESIZED_WIRE_80),
	.D33(SYNTHESIZED_WIRE_82),
	.D34(SYNTHESIZED_WIRE_1),
	.D35(SYNTHESIZED_WIRE_45),
	.D36(SYNTHESIZED_WIRE_61),
	.D37(SYNTHESIZED_WIRE_102),
	.D38(SYNTHESIZED_WIRE_57),
	.D39(SYNTHESIZED_WIRE_65),
	.D40(SYNTHESIZED_WIRE_94),
	.D41(SYNTHESIZED_WIRE_58),
	.D42(SYNTHESIZED_WIRE_83),
	.D43(SYNTHESIZED_WIRE_78),
	.D44(SYNTHESIZED_WIRE_66),
	.D45(SYNTHESIZED_WIRE_95),
	.D46(SYNTHESIZED_WIRE_103),
	.D47(SYNTHESIZED_WIRE_62),
	.D48(SYNTHESIZED_WIRE_86),
	.D49(SYNTHESIZED_WIRE_74),
	.D50(SYNTHESIZED_WIRE_90),
	.D51(SYNTHESIZED_WIRE_49),
	.D52(SYNTHESIZED_WIRE_46),
	.D53(SYNTHESIZED_WIRE_2),
	.D54(SYNTHESIZED_WIRE_53),
	.D55(SYNTHESIZED_WIRE_87),
	.D56(SYNTHESIZED_WIRE_75),
	.D57(SYNTHESIZED_WIRE_54),
	.D58(SYNTHESIZED_WIRE_69),
	.D59(SYNTHESIZED_WIRE_98),
	.D60(SYNTHESIZED_WIRE_50),
	.D61(SYNTHESIZED_WIRE_91),
	.D62(SYNTHESIZED_WIRE_79),
	.D63(SYNTHESIZED_WIRE_70),
	.D64(SYNTHESIZED_WIRE_99));

assign	SYNTHESIZED_WIRE_7 = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1 | SYNTHESIZED_WIRE_2 | SYNTHESIZED_WIRE_3;


rom_0111	b2v_inst10(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_4),
	.rom_out(SYNTHESIZED_WIRE_22));


rom_0110	b2v_inst11(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_5),
	.rom_out(SYNTHESIZED_WIRE_21));


rom_0101	b2v_inst12(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_6),
	.rom_out(SYNTHESIZED_WIRE_20));


rom_0100	b2v_inst13(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_7),
	.rom_out(SYNTHESIZED_WIRE_19));


rom_0011	b2v_inst14(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_8),
	.rom_out(SYNTHESIZED_WIRE_18));


rom_0010	b2v_inst15(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_9),
	.rom_out(SYNTHESIZED_WIRE_17));


rom_0001	b2v_inst16(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_10),
	.rom_out(SYNTHESIZED_WIRE_13));


rom_0000	b2v_inst17(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_11),
	.rom_out(SYNTHESIZED_WIRE_12));


or4bit	b2v_inst18(
	.in1(SYNTHESIZED_WIRE_12),
	.in2(SYNTHESIZED_WIRE_13),
	.out(SYNTHESIZED_WIRE_14));


or4bit	b2v_inst19(
	.in1(SYNTHESIZED_WIRE_14),
	.in2(SYNTHESIZED_WIRE_15),
	.out(SYNTHESIZED_WIRE_38));


rom_1111	b2v_inst2(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_16),
	.rom_out(SYNTHESIZED_WIRE_30));


or4bit	b2v_inst20(
	.in1(SYNTHESIZED_WIRE_17),
	.in2(SYNTHESIZED_WIRE_18),
	.out(SYNTHESIZED_WIRE_15));


or4bit	b2v_inst21(
	.in1(SYNTHESIZED_WIRE_19),
	.in2(SYNTHESIZED_WIRE_20),
	.out(SYNTHESIZED_WIRE_31));


or4bit	b2v_inst22(
	.in1(SYNTHESIZED_WIRE_21),
	.in2(SYNTHESIZED_WIRE_22),
	.out(SYNTHESIZED_WIRE_32));


or4bit	b2v_inst23(
	.in1(SYNTHESIZED_WIRE_23),
	.in2(SYNTHESIZED_WIRE_24),
	.out(SYNTHESIZED_WIRE_33));


or4bit	b2v_inst24(
	.in1(SYNTHESIZED_WIRE_25),
	.in2(SYNTHESIZED_WIRE_26),
	.out(SYNTHESIZED_WIRE_34));


or4bit	b2v_inst25(
	.in1(SYNTHESIZED_WIRE_27),
	.in2(SYNTHESIZED_WIRE_28),
	.out(SYNTHESIZED_WIRE_35));


or4bit	b2v_inst26(
	.in1(SYNTHESIZED_WIRE_29),
	.in2(SYNTHESIZED_WIRE_30),
	.out(SYNTHESIZED_WIRE_36));


or4bit	b2v_inst27(
	.in1(SYNTHESIZED_WIRE_31),
	.in2(SYNTHESIZED_WIRE_32),
	.out(SYNTHESIZED_WIRE_39));


or4bit	b2v_inst28(
	.in1(SYNTHESIZED_WIRE_33),
	.in2(SYNTHESIZED_WIRE_34),
	.out(SYNTHESIZED_WIRE_40));


or4bit	b2v_inst29(
	.in1(SYNTHESIZED_WIRE_35),
	.in2(SYNTHESIZED_WIRE_36),
	.out(SYNTHESIZED_WIRE_41));


rom_1110	b2v_inst3(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_37),
	.rom_out(SYNTHESIZED_WIRE_29));


or4bit	b2v_inst30(
	.in1(SYNTHESIZED_WIRE_38),
	.in2(SYNTHESIZED_WIRE_39),
	.out(SYNTHESIZED_WIRE_42));


or4bit	b2v_inst31(
	.in1(SYNTHESIZED_WIRE_40),
	.in2(SYNTHESIZED_WIRE_41),
	.out(SYNTHESIZED_WIRE_43));


or4bit	b2v_inst32(
	.in1(SYNTHESIZED_WIRE_42),
	.in2(SYNTHESIZED_WIRE_43),
	.out(sbox1_out));

assign	SYNTHESIZED_WIRE_37 = SYNTHESIZED_WIRE_44 | SYNTHESIZED_WIRE_45 | SYNTHESIZED_WIRE_46 | SYNTHESIZED_WIRE_47;

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_48 | SYNTHESIZED_WIRE_49 | SYNTHESIZED_WIRE_50 | SYNTHESIZED_WIRE_51;

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_52 | SYNTHESIZED_WIRE_53 | SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_55;

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57 | SYNTHESIZED_WIRE_58 | SYNTHESIZED_WIRE_59;

assign	SYNTHESIZED_WIRE_8 = SYNTHESIZED_WIRE_60 | SYNTHESIZED_WIRE_61 | SYNTHESIZED_WIRE_62 | SYNTHESIZED_WIRE_63;

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_64 | SYNTHESIZED_WIRE_65 | SYNTHESIZED_WIRE_66 | SYNTHESIZED_WIRE_67;

assign	SYNTHESIZED_WIRE_5 = SYNTHESIZED_WIRE_68 | SYNTHESIZED_WIRE_69 | SYNTHESIZED_WIRE_70 | SYNTHESIZED_WIRE_71;


rom_1101	b2v_inst4(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_72),
	.rom_out(SYNTHESIZED_WIRE_28));

assign	SYNTHESIZED_WIRE_4 = SYNTHESIZED_WIRE_73 | SYNTHESIZED_WIRE_74 | SYNTHESIZED_WIRE_75 | SYNTHESIZED_WIRE_76;

assign	SYNTHESIZED_WIRE_109 = SYNTHESIZED_WIRE_77 | SYNTHESIZED_WIRE_78 | SYNTHESIZED_WIRE_79 | SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_108 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_83 | SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_107 = SYNTHESIZED_WIRE_85 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_106 = SYNTHESIZED_WIRE_89 | SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_92;

assign	SYNTHESIZED_WIRE_105 = SYNTHESIZED_WIRE_93 | SYNTHESIZED_WIRE_94 | SYNTHESIZED_WIRE_95 | SYNTHESIZED_WIRE_96;

assign	SYNTHESIZED_WIRE_72 = SYNTHESIZED_WIRE_97 | SYNTHESIZED_WIRE_98 | SYNTHESIZED_WIRE_99 | SYNTHESIZED_WIRE_100;

assign	SYNTHESIZED_WIRE_16 = SYNTHESIZED_WIRE_101 | SYNTHESIZED_WIRE_102 | SYNTHESIZED_WIRE_103 | SYNTHESIZED_WIRE_104;


rom_1100	b2v_inst5(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_105),
	.rom_out(SYNTHESIZED_WIRE_27));


rom_1011	b2v_inst6(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_106),
	.rom_out(SYNTHESIZED_WIRE_26));


rom_1010	b2v_inst7(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_107),
	.rom_out(SYNTHESIZED_WIRE_25));


rom_1001	b2v_inst8(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_108),
	.rom_out(SYNTHESIZED_WIRE_24));


rom_1000	b2v_inst9(
	.clk(clk),
	.rst_n(rst_n),
	.sel(SYNTHESIZED_WIRE_109),
	.rom_out(SYNTHESIZED_WIRE_23));


endmodule
