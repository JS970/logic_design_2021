// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Nov 24 21:36:57 2021"

module Expension(
	e1,
	e2,
	e3,
	e4,
	e5,
	e6,
	e7,
	e8,
	e9,
	e10,
	e11,
	e12,
	e13,
	e14,
	e15,
	e16,
	e17,
	e18,
	e19,
	e20,
	e21,
	e22,
	e23,
	e24,
	e25,
	e26,
	e27,
	e28,
	e29,
	e30,
	e31,
	e32,
	eout1,
	eout2,
	eout3,
	eout4,
	eout5,
	eout6,
	eout7,
	eout8,
	eout9,
	eout10,
	eout11,
	eout12,
	eout13,
	eout14,
	eout15,
	eout16,
	eout17,
	eout18,
	eout19,
	eout20,
	eout21,
	eout22,
	eout23,
	eout24,
	eout25,
	eout26,
	eout27,
	eout28,
	eout29,
	eout30,
	eout31,
	eout32,
	eout33,
	eout34,
	eout35,
	eout36,
	eout37,
	eout38,
	eout39,
	eout40,
	eout41,
	eout42,
	eout43,
	eout44,
	eout45,
	eout46,
	eout47,
	eout48
);


input wire	e1;
input wire	e2;
input wire	e3;
input wire	e4;
input wire	e5;
input wire	e6;
input wire	e7;
input wire	e8;
input wire	e9;
input wire	e10;
input wire	e11;
input wire	e12;
input wire	e13;
input wire	e14;
input wire	e15;
input wire	e16;
input wire	e17;
input wire	e18;
input wire	e19;
input wire	e20;
input wire	e21;
input wire	e22;
input wire	e23;
input wire	e24;
input wire	e25;
input wire	e26;
input wire	e27;
input wire	e28;
input wire	e29;
input wire	e30;
input wire	e31;
input wire	e32;
output wire	eout1;
output wire	eout2;
output wire	eout3;
output wire	eout4;
output wire	eout5;
output wire	eout6;
output wire	eout7;
output wire	eout8;
output wire	eout9;
output wire	eout10;
output wire	eout11;
output wire	eout12;
output wire	eout13;
output wire	eout14;
output wire	eout15;
output wire	eout16;
output wire	eout17;
output wire	eout18;
output wire	eout19;
output wire	eout20;
output wire	eout21;
output wire	eout22;
output wire	eout23;
output wire	eout24;
output wire	eout25;
output wire	eout26;
output wire	eout27;
output wire	eout28;
output wire	eout29;
output wire	eout30;
output wire	eout31;
output wire	eout32;
output wire	eout33;
output wire	eout34;
output wire	eout35;
output wire	eout36;
output wire	eout37;
output wire	eout38;
output wire	eout39;
output wire	eout40;
output wire	eout41;
output wire	eout42;
output wire	eout43;
output wire	eout44;
output wire	eout45;
output wire	eout46;
output wire	eout47;
output wire	eout48;


assign	eout1 = e32;
assign	eout2 = e1;
assign	eout3 = e2;
assign	eout4 = e3;
assign	eout5 = e4;
assign	eout6 = e5;
assign	eout7 = e4;
assign	eout8 = e5;
assign	eout9 = e6;
assign	eout10 = e7;
assign	eout11 = e8;
assign	eout12 = e9;
assign	eout13 = e8;
assign	eout14 = e9;
assign	eout15 = e10;
assign	eout16 = e11;
assign	eout17 = e12;
assign	eout18 = e13;
assign	eout19 = e12;
assign	eout20 = e13;
assign	eout21 = e14;
assign	eout22 = e15;
assign	eout23 = e16;
assign	eout24 = e17;
assign	eout25 = e16;
assign	eout26 = e17;
assign	eout27 = e18;
assign	eout28 = e19;
assign	eout29 = e20;
assign	eout30 = e21;
assign	eout31 = e20;
assign	eout32 = e21;
assign	eout33 = e22;
assign	eout34 = e23;
assign	eout35 = e24;
assign	eout36 = e25;
assign	eout37 = e24;
assign	eout38 = e25;
assign	eout39 = e26;
assign	eout40 = e27;
assign	eout41 = e28;
assign	eout42 = e29;
assign	eout43 = e28;
assign	eout44 = e29;
assign	eout45 = e30;
assign	eout46 = e31;
assign	eout47 = e32;
assign	eout48 = e1;




endmodule
