// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Nov 24 20:56:12 2021"

module PC_2(
	pin1,
	pin2,
	pin3,
	pin4,
	pin5,
	pin6,
	pin7,
	pin8,
	pin9,
	pin10,
	pin11,
	pin12,
	pin13,
	pin14,
	pin15,
	pin16,
	pin17,
	pin18,
	pin19,
	pin20,
	pin21,
	pin22,
	pin23,
	pin24,
	pin25,
	pin26,
	pin27,
	pin28,
	pin29,
	pin30,
	pin31,
	pin32,
	pin33,
	pin34,
	pin35,
	pin36,
	pin37,
	pin38,
	pin39,
	pin40,
	pin41,
	pin42,
	pin43,
	pin44,
	pin45,
	pin46,
	pin47,
	pin48,
	pin49,
	pin50,
	pin51,
	pin52,
	pin53,
	pin54,
	pin55,
	pin56,
	pout1,
	pout2,
	pout3,
	pout4,
	pout5,
	pout6,
	pout7,
	pout8,
	pout9,
	pout10,
	pout11,
	pout12,
	pout13,
	pout14,
	pout15,
	pout16,
	pout17,
	pout18,
	pout19,
	pout20,
	pout21,
	pout22,
	pout23,
	pout24,
	pout25,
	pout26,
	pout27,
	pout28,
	pout29,
	pout30,
	pout31,
	pout32,
	pout33,
	pout34,
	pout35,
	pout36,
	pout37,
	pout38,
	pout39,
	pout40,
	pout41,
	pout42,
	pout43,
	pout44,
	pout45,
	pout46,
	pout47,
	pout48
);


input wire	pin1;
input wire	pin2;
input wire	pin3;
input wire	pin4;
input wire	pin5;
input wire	pin6;
input wire	pin7;
input wire	pin8;
input wire	pin9;
input wire	pin10;
input wire	pin11;
input wire	pin12;
input wire	pin13;
input wire	pin14;
input wire	pin15;
input wire	pin16;
input wire	pin17;
input wire	pin18;
input wire	pin19;
input wire	pin20;
input wire	pin21;
input wire	pin22;
input wire	pin23;
input wire	pin24;
input wire	pin25;
input wire	pin26;
input wire	pin27;
input wire	pin28;
input wire	pin29;
input wire	pin30;
input wire	pin31;
input wire	pin32;
input wire	pin33;
input wire	pin34;
input wire	pin35;
input wire	pin36;
input wire	pin37;
input wire	pin38;
input wire	pin39;
input wire	pin40;
input wire	pin41;
input wire	pin42;
input wire	pin43;
input wire	pin44;
input wire	pin45;
input wire	pin46;
input wire	pin47;
input wire	pin48;
input wire	pin49;
input wire	pin50;
input wire	pin51;
input wire	pin52;
input wire	pin53;
input wire	pin54;
input wire	pin55;
input wire	pin56;
output wire	pout1;
output wire	pout2;
output wire	pout3;
output wire	pout4;
output wire	pout5;
output wire	pout6;
output wire	pout7;
output wire	pout8;
output wire	pout9;
output wire	pout10;
output wire	pout11;
output wire	pout12;
output wire	pout13;
output wire	pout14;
output wire	pout15;
output wire	pout16;
output wire	pout17;
output wire	pout18;
output wire	pout19;
output wire	pout20;
output wire	pout21;
output wire	pout22;
output wire	pout23;
output wire	pout24;
output wire	pout25;
output wire	pout26;
output wire	pout27;
output wire	pout28;
output wire	pout29;
output wire	pout30;
output wire	pout31;
output wire	pout32;
output wire	pout33;
output wire	pout34;
output wire	pout35;
output wire	pout36;
output wire	pout37;
output wire	pout38;
output wire	pout39;
output wire	pout40;
output wire	pout41;
output wire	pout42;
output wire	pout43;
output wire	pout44;
output wire	pout45;
output wire	pout46;
output wire	pout47;
output wire	pout48;


assign	pout1 = pin14;
assign	pout2 = pin17;
assign	pout3 = pin11;
assign	pout4 = pin24;
assign	pout5 = pin1;
assign	pout6 = pin5;
assign	pout7 = pin3;
assign	pout8 = pin28;
assign	pout9 = pin15;
assign	pout10 = pin6;
assign	pout11 = pin21;
assign	pout12 = pin10;
assign	pout13 = pin23;
assign	pout14 = pin19;
assign	pout15 = pin12;
assign	pout16 = pin4;
assign	pout17 = pin26;
assign	pout18 = pin8;
assign	pout19 = pin16;
assign	pout20 = pin7;
assign	pout21 = pin27;
assign	pout22 = pin20;
assign	pout23 = pin13;
assign	pout24 = pin2;
assign	pout25 = pin41;
assign	pout26 = pin52;
assign	pout27 = pin31;
assign	pout28 = pin37;
assign	pout29 = pin47;
assign	pout30 = pin55;
assign	pout31 = pin30;
assign	pout32 = pin40;
assign	pout33 = pin51;
assign	pout34 = pin45;
assign	pout35 = pin33;
assign	pout36 = pin48;
assign	pout37 = pin44;
assign	pout38 = pin49;
assign	pout39 = pin39;
assign	pout40 = pin56;
assign	pout41 = pin34;
assign	pout42 = pin53;
assign	pout43 = pin46;
assign	pout44 = pin42;
assign	pout45 = pin50;
assign	pout46 = pin36;
assign	pout47 = pin29;
assign	pout48 = pin32;




endmodule
